#Software: 1.4.5 (commit 251f983)
#Command: breakdancer-max ZS97.bam.cfg 
#Library Statistics:
#/public07/yaowen/intansv/zs97_ncgr/ZS97.bam	mean:182.85	std:24.43	uppercutoff:261.07	lowercutoff:65.41	readlen:40	library:ZS97	reflen:375078573	seqcov:5.26656	phycov:12.0374	1:32040	2:206322	3:183193	4:15786	8:32442	32:97116
#Chr1	Pos1	Orientation1	Chr2	Pos2	Orientation2	Type	Size	Score	num_Reads	num_Reads_lib	ZS97.bam
chr05	65575	5+0-	chr05	65949	0+5-	DEL	353	88	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.04
chr05	86452	20+0-	chr05	87419	0+20-	DEL	988	99	20	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|20	NA
chr05	120264	7+2-	chr05	127693	6+6-	DEL	7382	83	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	1.07
chr05	120636	7+0-	chr05	120788	0+12-	DEL	95	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	0.16
chr05	153666	4+1-	chr05	153829	0+4-	DEL	107	80	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	1.84
chr05	197339	7+1-	chr05	197436	0+5-	DEL	99	93	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.23
chr05	201845	22+0-	chr05	201959	2+23-	DEL	114	99	22	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|22	0.20
chr05	208214	9+0-	chr05	208577	0+10-	DEL	354	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	0.11
chr05	226804	3+0-	chr05	226913	0+3-	DEL	86	55	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	1.69
chr05	230521	11+1-	chr05	230654	0+11-	DEL	136	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	0.18
chr05	276048	29+0-	chr05	276182	0+29-	DEL	148	99	29	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|29	0.45
chr05	276751	2+0-	chr05	276950	0+2-	DEL	137	47	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	1.30
chr05	280404	8+0-	chr05	281218	0+7-	DEL	739	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	0.13
chr05	334347	5+0-	chr05	334632	0+5-	DEL	285	86	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.05
chr05	340558	3+1-	chr05	347164	0+2-	DEL	6593	45	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	2.61
chr05	348417	13+0-	chr05	350116	0+13-	DEL	1683	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	0.04
chr05	366435	14+0-	chr05	367950	0+14-	DEL	1521	99	14	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|14	0.02
chr05	379192	25+0-	chr05	404522	0+25-	DEL	25322	99	25	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|25	NA
chr05	405042	11+0-	chr05	408729	0+11-	DEL	3689	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	NA
chr05	470271	5+5-	chr05	470628	5+5-	DEL	85	69	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	NA
chr05	484719	24+0-	chr05	484861	0+24-	DEL	138	99	24	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|24	0.26
chr05	498607	14+0-	chr05	505453	0+14-	DEL	6832	99	14	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|14	0.26
chr05	541621	7+0-	chr05	541721	6+6-	DEL	95	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.11
chr05	541807	6+6-	chr05	542031	0+7-	DEL	201	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.23
chr05	582645	3+0-	chr05	582811	0+3-	DEL	123	60	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.60
chr05	614084	16+0-	chr05	628895	2+16-	DEL	14846	99	16	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|16	NA
chr05	657418	4+1-	chr05	657497	0+3-	DEL	88	50	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	2.27
chr05	664197	2+0-	chr05	664346	1+2-	DEL	81	51	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	2.31
chr05	665958	12+0-	chr05	667136	0+12-	DEL	1196	99	12	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|12	NA
chr05	681547	5+0-	chr05	683014	0+5-	DEL	1441	90	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.03
chr05	700037	5+0-	chr05	700312	0+5-	DEL	218	97	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	NA
chr05	706435	11+0-	chr05	707841	0+11-	DEL	1399	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	0.04
chr05	822333	3+0-	chr05	822437	0+3-	DEL	86	54	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	1.09
chr05	861533	0+4-	chr05	861582	0+4-	INV	-99	72	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	915043	2+0-	chr05	917776	0+2-	DEL	2644	57	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.04
chr05	972863	10+0-	chr05	977659	0+10-	DEL	4796	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	12.52
chr05	974945	1+4-	chr05	975011	1+4-	INV	-105	70	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	1009748	2+0-	chr05	1009875	1+2-	DEL	90	47	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	1.22
chr05	1091289	5+0-	chr05	1102799	0+5-	DEL	11484	91	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.00
chr05	1112010	4+0-	chr05	1112183	0+4-	DEL	95	98	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	1.75
chr05	1115271	3+0-	chr05	1115408	2+5-	DEL	89	51	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	2.21
chr05	1152575	3+0-	chr05	1152712	0+3-	DEL	90	61	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	1.68
chr05	1155009	21+0-	chr05	1155565	0+21-	DEL	561	99	21	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|21	0.05
chr05	1161457	4+2-	chr05	1161609	0+4-	DEL	91	86	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	2.11
chr05	1166830	6+0-	chr05	1168062	0+6-	DEL	1160	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.08
chr05	1291603	0+6-	chr05	1291649	0+6-	INV	-105	99	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	NA
chr05	1302899	18+0-	chr05	1305821	0+18-	DEL	2910	99	18	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|18	0.03
chr05	1386815	16+0-	chr05	1389331	0+16-	DEL	2519	99	16	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|16	0.02
chr05	1409610	25+0-	chr05	1412844	0+25-	DEL	3245	99	25	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|25	0.01
chr05	1442743	16+0-	chr05	1443102	0+16-	DEL	326	99	16	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|16	0.23
chr05	1464922	7+0-	chr05	1465219	0+7-	DEL	284	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	0.05
chr05	1491177	28+0-	chr05	1491595	0+27-	DEL	442	99	27	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|27	NA
chr05	1530688	13+0-	chr05	1530829	0+13-	DEL	142	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	0.09
chr05	1685654	9+0-	chr05	1686167	0+9-	DEL	505	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	0.03
chr05	1688921	21+0-	chr05	1696567	4+21-	DEL	7664	99	21	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|21	NA
chr05	1709745	10+0-	chr05	1709978	18+10-	DEL	184	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	0.57
chr05	1710156	18+10-	chr05	1710425	0+18-	DEL	268	99	18	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|18	NA
chr05	1712267	4+0-	chr05	1712538	0+4-	DEL	234	78	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.05
chr05	1733342	3+0-	chr05	1733578	0+3-	DEL	158	75	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.45
chr05	1766811	18+0-	chr05	1778172	0+18-	DEL	11345	99	18	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|18	NA
chr05	1783486	11+0-	chr05	1784891	0+11-	DEL	1375	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	0.01
chr05	1797984	13+0-	chr05	1802325	0+13-	DEL	4341	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	0.01
chr05	1802845	22+0-	chr05	1803476	0+22-	DEL	633	99	22	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|22	0.14
chr05	1809475	3+0-	chr05	1809938	0+3-	DEL	374	82	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.03
chr05	1828254	6+0-	chr05	1828406	0+6-	DEL	141	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	NA
chr05	1839141	8+0-	chr05	1839749	0+8-	DEL	524	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.05
chr05	1921493	8+0-	chr05	1922917	0+8-	DEL	1413	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.05
chr05	2019472	17+0-	chr05	2019716	0+17-	DEL	238	99	17	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|17	NA
chr05	2020503	2+0-	chr05	2020806	1+2-	DEL	232	55	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	2030039	2+0-	chr05	2030383	0+2-	DEL	279	47	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.28
chr05	2032386	15+0-	chr05	2044616	0+15-	DEL	12225	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	0.00
chr05	2049414	7+0-	chr05	2049880	0+7-	DEL	451	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	0.06
chr05	2076230	7+0-	chr05	2076538	0+7-	DEL	299	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	0.13
chr05	2081872	3+0-	chr05	2081961	2+3-	DEL	99	48	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.12
chr05	2094543	4+1-	chr05	2094669	2+3-	DEL	91	44	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	2.36
chr05	2112637	2+0-	chr05	2112808	2+3-	DEL	87	53	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	1.77
chr05	2119684	24+1-	chr05	2119838	0+24-	DEL	147	99	24	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|24	0.08
chr05	2120425	3+0-	chr05	2120815	0+3-	DEL	310	75	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.36
chr05	2121948	6+0-	chr05	2122082	0+6-	DEL	105	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.09
chr05	2123832	9+0-	chr05	2128080	1+9-	DEL	4248	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	0.01
chr05	2131355	9+0-	chr05	2133569	0+13-	DEL	2153	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	NA
chr05	2232719	16+0-	chr05	2239174	0+16-	DEL	6457	99	16	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|16	NA
chr05	2248980	12+12-	chr05	2249334	12+12-	DEL	94	99	12	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|12	NA
chr05	2270521	13+1-	chr05	2283410	0+13-	DEL	12884	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	NA
chr05	2298634	8+0-	chr05	2299026	0+8-	DEL	337	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.21
chr05	2308966	8+0-	chr05	2309128	0+8-	DEL	157	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.08
chr05	2321120	2+0-	chr05	2321860	2+4-	DEL	664	54	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.14
chr05	2328591	13+0-	chr05	2328719	0+12-	DEL	168	99	12	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|12	NA
chr05	2362216	15+0-	chr05	2362472	1+16-	DEL	231	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	NA
chr05	2405013	6+0-	chr05	2416431	0+6-	DEL	11338	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	NA
chr05	2437971	5+0-	chr05	2439220	0+5-	DEL	1192	99	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.01
chr05	2453626	23+0-	chr05	2460061	0+23-	DEL	6435	99	23	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|23	0.00
chr05	2472976	22+0-	chr05	2477807	0+22-	DEL	4841	99	22	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|22	0.00
chr05	2485527	5+0-	chr05	2485632	3+5-	DEL	85	90	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	1.19
chr05	2562923	0+2-	chr05	2563067	0+2-	INV	-42	82	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	2.29
chr05	2567373	7+0-	chr05	2567532	0+7-	DEL	98	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	0.70
chr05	2584226	4+0-	chr05	2584259	4+0-	INV	-114	75	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	2594055	3+2-	chr05	2594290	0+3-	DEL	150	62	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.06
chr05	2634491	10+0-	chr05	2634614	0+10-	DEL	94	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	0.87
chr05	2636234	13+7-	chr05	2637171	0+13-	DEL	1056	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	0.23
chr05	2678840	10+0-	chr05	2679344	0+10-	DEL	458	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	0.20
chr05	2686821	4+0-	chr05	2698636	0+4-	DEL	11767	76	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.00
chr05	2741220	15+1-	chr05	2741488	0+16-	DEL	221	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	0.20
chr05	2748901	15+0-	chr05	2753063	1+17-	DEL	4153	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	0.00
chr05	2754781	26+0-	chr05	2755040	0+26-	DEL	244	99	26	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|26	0.26
chr05	2755811	17+0-	chr05	2756134	0+17-	DEL	311	99	17	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|17	0.13
chr05	2758521	6+0-	chr05	2760125	0+5-	DEL	1567	93	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.02
chr05	2761545	17+1-	chr05	2762613	0+16-	DEL	1019	99	16	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|16	0.06
chr05	2797477	12+0-	chr05	2803733	0+12-	DEL	6246	99	12	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|12	NA
chr05	2808330	15+1-	chr05	2809386	0+15-	DEL	1095	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	NA
chr05	2867281	2+0-	chr05	2867477	2+0-	INV	-2	75	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	3.35
chr05	2890771	22+0-	chr05	2891012	0+22-	DEL	245	99	22	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|22	NA
chr05	2945387	15+0-	chr05	2952291	0+15-	DEL	6906	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	NA
chr05	2955552	7+1-	chr05	2964340	1+7-	DEL	8779	90	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.01
chr05	2982127	14+0-	chr05	2983579	0+14-	DEL	1461	99	14	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|14	0.01
chr05	2986916	15+0-	chr05	2987435	1+16-	DEL	503	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	0.08
chr05	2994956	6+0-	chr05	2995095	0+6-	DEL	127	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.35
chr05	2999151	8+1-	chr05	3003345	1+7-	DEL	4200	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	0.01
chr05	3008104	9+0-	chr05	3008231	0+9-	DEL	96	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	0.75
chr05	3016418	2+0-	chr05	3029744	0+2-	DEL	13234	59	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	3067944	6+0-	chr05	3068646	0+6-	DEL	673	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.19
chr05	3077399	3+0-	chr05	3077528	1+3-	DEL	89	54	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	1.20
chr05	3088652	6+0-	chr05	3088782	0+6-	DEL	94	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	1.66
chr05	3104311	4+0-	chr05	3104366	4+0-	INV	-92	71	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	3109159	19+0-	chr05	3109578	0+19-	DEL	426	99	19	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|19	0.13
chr05	3125229	18+0-	chr05	3125419	2+17-	DEL	163	99	17	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|17	0.47
chr05	3163532	20+0-	chr05	3163761	1+20-	DEL	263	99	20	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|20	0.06
chr05	3176843	6+0-	chr05	3176991	0+6-	DEL	83	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.75
chr05	3182222	0+4-	chr05	3182279	0+4-	INV	-90	71	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	3223779	3+0-	chr05	3229630	0+3-	DEL	5800	61	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	NA
chr05	3233358	3+0-	chr05	3233546	0+3-	DEL	144	59	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.48
chr05	3243936	19+1-	chr05	3244148	0+19-	DEL	263	99	19	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|19	0.43
chr05	3300982	10+2-	chr05	3301301	0+10-	DEL	310	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	0.13
chr05	3326524	6+0-	chr05	3326584	6+0-	INV	-87	97	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	NA
chr05	3335043	5+0-	chr05	3335426	0+6-	DEL	326	99	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	NA
chr05	3358702	8+0-	chr05	3358836	0+8-	DEL	93	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	1.26
chr05	3447479	16+0-	chr05	3447753	0+16-	DEL	280	99	16	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|16	0.05
chr05	3523209	4+0-	chr05	3523344	0+4-	DEL	82	83	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	1.97
chr05	3625428	5+1-	chr05	3626107	1+5-	DEL	792	73	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	NA
chr05	3668983	4+0-	chr05	3669204	4+0-	INV	-8	58	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	3783456	18+0-	chr05	3784609	17+19-	DEL	1307	99	18	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|18	0.08
chr05	3744052	10+0-	chr05	3751972	0+10-	DEL	7928	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	0.00
chr05	3774641	7+0-	chr05	3774736	0+7-	DEL	88	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	0.23
chr05	3777927	2+0-	chr05	3778005	3+4-	DEL	83	42	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	1.08
chr05	3778151	3+4-	chr05	3778229	0+3-	DEL	85	60	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	2.55
chr05	3791166	13+0-	chr05	3798249	0+13-	DEL	7090	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	NA
chr05	3810951	11+0-	chr05	3811207	0+11-	DEL	255	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	NA
chr05	3860406	20+1-	chr05	3867103	0+19-	DEL	6679	99	19	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|19	0.00
chr05	3882000	15+0-	chr05	3889940	9+13-	DEL	7952	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	NA
chr05	3882000	15+0-	chr05	3890294	0+11-	DEL	8194	35	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.00
chr05	3890060	9+13-	chr05	3890294	0+11-	DEL	213	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	0.06
chr05	3895046	4+0-	chr05	3931951	12+4-	DEL	36859	64	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.00
chr05	3932165	12+4-	chr05	3955351	1+14-	DEL	23192	99	12	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|12	0.00
chr05	3960111	5+0-	chr05	3964126	0+5-	DEL	4010	86	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.01
chr05	3965450	6+0-	chr05	3965677	0+6-	DEL	145	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.06
chr05	4033770	13+0-	chr05	4045044	1+13-	DEL	11303	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	0.00
chr05	4074846	13+0-	chr05	4076032	2+13-	DEL	1158	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	1.01
chr05	4076204	2+13-	chr05	4076354	0+2-	DEL	102	37	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	5.58
chr05	4089795	4+0-	chr05	4089958	0+3-	DEL	84	74	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.38
chr05	4368561	2+0-	chr05	4370796	24+2-	DEL	2402	32	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	5.84
chr05	4135661	12+0-	chr05	4136019	0+12-	DEL	343	99	12	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|12	NA
chr05	4151856	21+0-	chr05	4152294	0+21-	DEL	447	99	21	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|21	NA
chr05	4155922	3+0-	chr05	4156695	0+3-	DEL	681	84	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	NA
chr05	4178028	8+0-	chr05	4178551	1+9-	DEL	465	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.08
chr05	4187967	6+0-	chr05	4188351	0+6-	DEL	354	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	NA
chr05	4194682	5+0-	chr05	4195025	0+6-	DEL	318	87	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.08
chr05	4250987	14+0-	chr05	4253130	0+14-	DEL	2133	99	14	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|14	0.02
chr05	4255220	5+1-	chr05	4255390	5+1-	INV	-113	60	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	4275555	16+1-	chr05	4278733	1+16-	DEL	3253	99	16	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|16	NA
chr05	4333064	13+0-	chr05	4344215	0+13-	DEL	11131	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	0.00
chr05	4353765	7+0-	chr05	4356935	0+6-	DEL	3151	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.00
chr05	4369252	14+0-	chr05	4369687	2+13-	DEL	471	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	3.49
chr05	4396018	3+0-	chr05	4401859	0+3-	DEL	5783	61	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.01
chr05	4409514	7+0-	chr05	4410685	0+7-	DEL	1101	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	0.04
chr05	4432415	11+0-	chr05	4435568	0+11-	DEL	3140	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	0.00
chr05	4479498	17+2-	chr05	4479586	0+17-	DEL	95	99	17	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|17	0.74
chr05	4551622	5+1-	chr05	4552298	0+5-	DEL	626	99	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.09
chr05	4598787	6+0-	chr05	4599694	0+6-	DEL	839	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	NA
chr05	4636331	20+0-	chr05	4644051	0+20-	DEL	7714	99	20	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|20	0.01
chr05	4686908	4+0-	chr05	4686983	2+4-	DEL	89	66	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	1.66
chr05	4712000	17+0-	chr05	4712621	0+17-	DEL	631	99	17	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|17	0.05
chr05	4870141	4+0-	chr05	4870205	4+0-	INV	-83	70	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	4925179	9+0-	chr05	4925837	2+10-	DEL	696	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	1.64
chr05	5224539	2+0-	chr05	5225232	2+0-	INV	505	79	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	2.34
chr05	5307544	2+0-	chr05	5307777	2+0-	INV	19	66	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	2.55
chr05	5404454	3+0-	chr05	5410038	1+7-	DEL	5495	64	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	NA
chr05	5405132	4+0-	chr05	5410038	1+7-	DEL	4868	84	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	NA
chr05	5446036	11+0-	chr05	5446160	0+11-	DEL	95	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	0.67
chr05	5550261	0+16-	chr05	5550392	0+16-	INV	-52	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	NA
chr05	5555551	22+0-	chr05	5557245	0+22-	DEL	1699	99	22	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|22	NA
chr05	5622270	5+0-	chr05	5646085	0+5-	DEL	23795	89	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.00
chr05	5660955	8+0-	chr05	5671854	0+8-	DEL	10879	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.00
chr05	5698786	10+1-	chr05	5698934	0+10-	DEL	109	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	0.91
chr05	5850682	5+0-	chr05	5851835	0+5-	DEL	1116	97	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.06
chr05	6001735	8+0-	chr05	6002058	0+8-	DEL	249	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.25
chr05	6013417	4+0-	chr05	6014345	0+4-	DEL	847	98	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.17
chr05	6033137	18+0-	chr05	6040489	0+18-	DEL	7356	99	18	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|18	0.02
chr05	6052582	8+0-	chr05	6052946	0+8-	DEL	332	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.04
chr05	6104849	5+0-	chr05	6104927	0+5-	DEL	88	82	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.27
chr05	6105948	13+0-	chr05	6106913	0+13-	DEL	984	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	NA
chr05	6139630	16+0-	chr05	6140223	0+16-	DEL	595	99	16	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|16	NA
chr05	6169799	10+0-	chr05	6170314	0+8-	DEL	493	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.03
chr05	6172147	3+0-	chr05	6172787	2+3-	DEL	567	71	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.07
chr05	6195004	5+0-	chr05	6195311	0+5-	DEL	283	86	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.09
chr05	6197871	7+1-	chr05	6203200	0+7-	DEL	5346	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	0.02
chr05	6212735	4+2-	chr05	6212912	0+4-	DEL	95	69	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.29
chr05	6299975	13+0-	chr05	6300119	1+14-	DEL	119	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	0.17
chr05	6323348	8+0-	chr05	6324003	0+9-	DEL	646	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.04
chr05	6327038	7+0-	chr05	6327174	1+8-	DEL	90	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	1.24
chr05	6329115	4+0-	chr05	6329177	4+0-	INV	-85	70	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	6394381	15+0-	chr05	6395366	0+15-	DEL	974	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	0.04
chr05	6470908	0+4-	chr05	6470937	0+4-	INV	-154	86	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	6477593	0+4-	chr05	6477659	0+4-	INV	-81	70	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	6646319	0+6-	chr05	6646404	0+6-	INV	-66	67	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	6691561	4+0-	chr05	6691600	4+0-	INV	-108	74	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	6747900	10+0-	chr05	6748030	0+10-	DEL	124	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	0.28
chr05	6764484	4+0-	chr05	6765086	1+5-	DEL	518	91	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.21
chr05	6765540	2+0-	chr05	6765660	0+2-	DEL	81	41	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.59
chr05	6770164	23+1-	chr05	6773110	0+23-	DEL	2982	99	23	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|23	NA
chr05	6818932	18+2-	chr05	6819130	0+17-	DEL	189	99	17	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|17	0.39
chr05	6827063	2+0-	chr05	6827158	0+3-	DEL	84	37	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	2.92
chr05	6841431	7+0-	chr05	6841672	1+7-	DEL	256	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	0.39
chr05	6845893	20+0-	chr05	6846051	0+20-	DEL	155	99	20	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|20	0.24
chr05	6852355	3+0-	chr05	6852554	0+3-	DEL	102	90	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.52
chr05	6872252	2+0-	chr05	6874614	0+2-	DEL	2272	59	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	6880235	6+0-	chr05	6880451	2+6-	DEL	149	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.61
chr05	6880530	2+6-	chr05	6881048	3+2-	DEL	414	37	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.08
chr05	6910121	9+1-	chr05	6913128	7+9-	DEL	2984	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	NA
chr05	6913325	7+9-	chr05	6913921	0+7-	DEL	593	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	NA
chr05	6942362	5+0-	chr05	6944726	5+0-	INV	2186	99	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	1.01
chr05	6949299	11+0-	chr05	6949776	0+11-	DEL	469	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	0.12
chr05	6953793	6+0-	chr05	6954018	0+6-	DEL	158	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	1.05
chr05	6960074	7+2-	chr05	6960183	0+5-	DEL	89	77	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	1.90
chr05	6963161	6+0-	chr05	6963357	0+6-	DEL	125	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.07
chr05	7018668	8+1-	chr05	7019214	1+7-	DEL	511	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	NA
chr05	7028787	11+0-	chr05	7029013	0+11-	DEL	242	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	NA
chr05	7061829	10+0-	chr05	7061989	0+10-	DEL	167	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	NA
chr05	7114320	16+0-	chr05	7114715	0+16-	DEL	371	99	16	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|16	0.14
chr05	7122590	4+0-	chr05	7122683	0+4-	DEL	103	65	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.71
chr05	7182462	9+0-	chr05	7187757	1+10-	DEL	5246	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	0.01
chr05	7236237	4+0-	chr05	7236400	0+4-	DEL	92	49	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.61
chr05	7259663	3+0-	chr05	7266413	0+3-	DEL	6692	64	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.00
chr05	7300248	8+0-	chr05	7300342	0+9-	DEL	118	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.12
chr05	7394062	2+1-	chr05	7394373	0+2-	DEL	228	54	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.26
chr05	7539257	12+0-	chr05	7550284	0+12-	DEL	11011	99	12	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|12	0.00
chr05	7550570	0+4-	chr05	7550628	0+4-	INV	-89	71	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	7556935	9+0-	chr05	7557284	0+9-	DEL	358	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	NA
chr05	7626573	13+0-	chr05	7627051	11+13-	DEL	469	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	0.03
chr05	7627213	11+13-	chr05	7627953	0+11-	DEL	719	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	0.02
chr05	7657548	3+3-	chr05	7657594	3+3-	INV	-142	72	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	7719567	9+0-	chr05	7719864	0+9-	DEL	255	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	0.23
chr05	7753048	4+0-	chr05	7753141	0+3-	DEL	91	61	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.83
chr05	7787302	9+0-	chr05	7798420	0+9-	DEL	11115	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	0.01
chr05	7818983	11+7-	chr05	7819270	9+8-	DEL	355	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	NA
chr05	7819373	9+8-	chr05	7819713	0+10-	DEL	331	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	NA
chr05	8042923	8+0-	chr05	8043423	0+6-	DEL	486	66	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.11
chr05	7862090	19+0-	chr05	7862235	0+19-	DEL	138	99	19	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|19	0.51
chr05	7865041	16+1-	chr05	7865293	1+16-	DEL	250	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	0.05
chr05	7879404	3+0-	chr05	7879592	0+3-	DEL	101	74	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.07
chr05	7975861	13+0-	chr05	7975970	1+13-	DEL	99	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	0.63
chr05	7979557	13+0-	chr05	7979826	1+13-	DEL	259	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	0.10
chr05	7980481	11+0-	chr05	7980691	0+11-	DEL	210	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	NA
chr05	7997604	18+0-	chr05	7997849	0+18-	DEL	232	99	18	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|18	0.33
chr05	8007921	13+0-	chr05	8008901	0+13-	DEL	977	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	0.04
chr05	8010226	19+0-	chr05	8010465	1+21-	DEL	237	99	19	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|19	NA
chr05	8026040	12+1-	chr05	8026229	0+11-	DEL	106	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	0.07
chr05	8027076	9+0-	chr05	8027707	0+8-	DEL	607	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	NA
chr05	8053367	9+0-	chr05	8057264	0+8-	DEL	3832	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.01
chr05	8064856	4+1-	chr05	8077886	0+3-	DEL	12957	56	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	NA
chr05	8086492	4+0-	chr05	8086513	4+0-	INV	-126	77	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	8107256	3+0-	chr05	8107366	0+3-	DEL	86	55	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	1.68
chr05	8134253	0+2-	chr05	8135835	0+2-	INV	1402	85	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.04
chr05	8159764	10+0-	chr05	8171552	0+11-	DEL	11756	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	0.01
chr05	8174953	12+0-	chr05	8175614	0+13-	DEL	603	99	12	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|12	NA
chr05	8189772	20+0-	chr05	8189973	0+20-	DEL	182	99	20	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|20	0.06
chr05	8198731	0+2-	chr05	8199559	0+2-	INV	652	72	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	1.76
chr05	8223572	5+0-	chr05	8223691	0+4-	DEL	83	65	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	1.58
chr05	8255960	22+0-	chr05	8259900	8+22-	DEL	3929	99	22	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|22	0.01
chr05	8260207	8+22-	chr05	8260760	0+8-	DEL	498	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	NA
chr05	8297710	20+0-	chr05	8298371	0+20-	DEL	660	99	20	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|20	NA
chr05	8354013	2+0-	chr05	8354149	2+0-	INV	-11	69	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	1.07
chr05	8394367	17+2-	chr05	8394757	1+16-	DEL	493	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	0.61
chr05	8395491	12+0-	chr05	8396032	0+12-	DEL	518	99	12	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|12	1.16
chr05	8488196	4+0-	chr05	8488252	4+0-	INV	-91	71	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	8535231	18+0-	chr05	8535343	0+19-	DEL	118	99	18	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|18	0.10
chr05	8560033	14+0-	chr05	8563664	2+16-	DEL	3622	99	14	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|14	0.01
chr05	8580267	4+0-	chr05	8580669	0+4-	DEL	311	99	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.10
chr05	8665869	3+0-	chr05	8670166	0+3-	DEL	4264	57	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	NA
chr05	8696879	7+0-	chr05	8697513	0+8-	DEL	582	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	0.02
chr05	8701290	1+3-	chr05	8702396	1+3-	INV	936	56	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	1.41
chr05	8702150	2+0-	chr05	8702230	1+3-	DEL	90	40	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.40
chr05	8717562	8+0-	chr05	8729838	0+8-	DEL	12218	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.01
chr05	8736157	15+0-	chr05	8748114	0+14-	DEL	11923	99	14	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|14	0.01
chr05	8759307	8+0-	chr05	8766832	0+8-	DEL	7444	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	NA
chr05	8789753	3+0-	chr05	8838116	0+3-	DEL	48293	67	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.00
chr05	8894909	17+0-	chr05	8898059	0+17-	DEL	3134	99	17	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|17	0.00
chr05	8921400	24+1-	chr05	8927803	0+23-	DEL	6413	99	23	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|23	0.01
chr05	8961020	12+0-	chr05	8962328	0+12-	DEL	1290	99	12	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|12	NA
chr05	8963166	2+6-	chr05	8963349	2+6-	INV	-134	60	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	10117263	2+0-	chr05	10117523	2+2-	INV	-32	86	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	1.34
chr05	10118349	2+2-	chr05	10118384	2+2-	INV	-182	83	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	10356312	4+0-	chr05	10356356	4+0-	INV	-103	73	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	10529330	1+4-	chr05	10529391	1+4-	INV	-86	70	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	3215974	3+2-	chr05	11733519	2+5-	DEL	8517499	60	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	1.77
chr05	11445411	6+0-	chr05	11445615	1+7-	DEL	209	93	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	2.80
chr05	11480921	2+0-	chr05	11481231	2+2-	INV	57	84	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	1.54
chr05	11974340	3+1-	chr05	11974626	3+1-	INV	-13	61	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	2.18
chr05	12014477	0+6-	chr05	12016019	0+6-	INV	1334	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	5.41
chr05	12886638	16+0-	chr05	12892009	0+16-	DEL	5367	99	16	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|16	NA
chr05	13089762	0+4-	chr05	13089811	0+4-	INV	-98	72	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	13142936	8+1-	chr05	13180473	0+8-	DEL	37506	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.03
chr05	13291698	0+8-	chr05	13291837	0+8-	INV	-35	87	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	NA
chr05	13644780	22+0-	chr05	13655489	4+20-	DEL	10703	99	20	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|20	0.00
chr05	13717366	0+4-	chr05	13717369	0+4-	INV	-144	82	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	13831875	0+4-	chr05	13831892	0+4-	INV	-130	78	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	13864304	5+0-	chr05	13864433	0+5-	DEL	140	84	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.09
chr05	14038691	5+0-	chr05	14038849	5+0-	INV	-134	61	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	14089207	17+0-	chr05	14100870	0+17-	DEL	11625	99	17	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|17	NA
chr05	14116903	22+0-	chr05	14129776	0+22-	DEL	12879	99	22	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|22	0.00
chr05	14255460	13+0-	chr05	14258839	0+13-	DEL	3363	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	0.00
chr05	14305803	9+0-	chr05	14306869	0+9-	DEL	1018	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	0.04
chr05	14310676	2+0-	chr05	14310858	0+2-	DEL	89	60	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	3.85
chr05	14358165	9+0-	chr05	14358236	0+9-	DEL	93	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	0.86
chr05	14746362	30+1-	chr05	14747195	0+30-	DEL	868	99	30	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|30	0.04
chr05	14748598	17+0-	chr05	14748856	0+17-	DEL	245	99	17	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|17	0.16
chr05	14759303	8+0-	chr05	14777629	0+8-	DEL	18301	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	NA
chr05	14813090	15+0-	chr05	14813205	0+15-	DEL	106	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	0.61
chr05	14877294	4+0-	chr05	14878000	0+4-	DEL	668	79	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	NA
chr05	14910155	6+0-	chr05	14910428	0+6-	DEL	271	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	NA
chr05	14920375	21+10-	chr05	14920486	0+10-	DEL	101	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	0.10
chr05	14933025	12+0-	chr05	14933894	0+12-	DEL	800	99	12	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|12	0.17
chr05	14944901	1+1-	chr05	14945177	2+2-	INV	1	66	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	1.32
chr05	14946900	14+0-	chr05	14947410	0+14-	DEL	485	99	14	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|14	0.11
chr05	14984813	9+0-	chr05	14985184	0+9-	DEL	352	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	0.26
chr05	14992058	7+0-	chr05	14992563	1+8-	DEL	505	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	NA
chr05	14999346	4+0-	chr05	14999368	4+0-	INV	-125	77	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	15034033	13+0-	chr05	15034127	2+15-	DEL	93	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	0.24
chr05	15092329	4+0-	chr05	15157598	4+0-	INV	65072	99	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	1.74
chr05	15125378	2+6-	chr05	15125468	2+6-	INV	-57	67	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	15146546	4+1-	chr05	15146728	4+1-	INV	-57	60	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	15166574	6+0-	chr05	15166647	0+6-	DEL	88	98	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.14
chr05	15254567	5+0-	chr05	15265162	1+4-	DEL	10527	95	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.00
chr05	15292483	3+0-	chr05	15305193	0+3-	DEL	12621	81	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.00
chr05	15472898	12+0-	chr05	15480744	0+12-	DEL	7839	99	12	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|12	0.00
chr05	15488673	6+0-	chr05	15488937	0+6-	DEL	237	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.20
chr05	15489995	22+1-	chr05	15491267	0+22-	DEL	1301	99	22	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|22	0.01
chr05	15544394	6+2-	chr05	15552128	0+7-	DEL	7722	63	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.00
chr05	15547820	3+1-	chr05	15552128	0+7-	DEL	4292	61	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.01
chr05	15577573	8+0-	chr05	15577679	1+9-	DEL	96	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.32
chr05	15604187	13+0-	chr05	15606484	0+13-	DEL	2260	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	0.04
chr05	15711137	11+0-	chr05	15722178	0+11-	DEL	10989	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	0.00
chr05	15741849	21+0-	chr05	15742203	0+21-	DEL	342	99	21	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|21	0.16
chr05	15744453	14+0-	chr05	15744663	0+14-	DEL	191	99	14	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|14	0.19
chr05	15755057	4+0-	chr05	15755080	4+0-	INV	-124	77	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	15774103	4+0-	chr05	15774373	0+4-	DEL	218	82	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	NA
chr05	15824859	19+0-	chr05	15828923	0+19-	DEL	4045	99	19	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|19	0.00
chr05	15844411	19+0-	chr05	15863727	0+19-	DEL	19319	99	19	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|19	0.00
chr05	15882438	0+4-	chr05	15882494	0+4-	INV	-91	71	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	15895353	21+0-	chr05	15895437	0+21-	DEL	98	99	21	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|21	0.38
chr05	15963088	2+0-	chr05	15977432	0+2-	DEL	14269	51	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.00
chr05	16004283	3+0-	chr05	16010925	1+4-	DEL	6630	49	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	NA
chr05	16023971	13+1-	chr05	16024346	0+12-	DEL	370	99	12	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|12	0.07
chr05	16029841	16+0-	chr05	16041095	15+16-	DEL	11241	99	16	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|16	0.00
chr05	16041315	15+16-	chr05	16041449	0+15-	DEL	141	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	NA
chr05	16060015	3+0-	chr05	16070459	0+3-	DEL	10426	55	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.01
chr05	16081695	6+0-	chr05	16081772	0+6-	DEL	90	98	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.68
chr05	16082244	14+0-	chr05	16083548	0+14-	DEL	1280	99	14	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|14	0.07
chr05	16086164	6+0-	chr05	16086306	0+6-	DEL	90	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	2.15
chr05	16086680	17+1-	chr05	16086811	0+16-	DEL	97	99	16	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|16	0.18
chr05	16248379	4+0-	chr05	16249218	0+5-	DEL	817	80	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.09
chr05	16276358	0+4-	chr05	16276409	0+4-	INV	-98	72	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	16343713	2+0-	chr05	16343812	1+3-	DEL	82	45	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	2.49
chr05	16376610	5+0-	chr05	16376949	0+5-	DEL	340	85	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.12
chr05	16399509	4+0-	chr05	16419850	0+4-	DEL	20279	90	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.01
chr05	16426421	4+0-	chr05	16431774	1+4-	DEL	5340	76	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.18
chr05	16433145	12+0-	chr05	16437333	0+12-	DEL	4198	99	12	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|12	NA
chr05	16464307	5+0-	chr05	16464490	0+5-	DEL	95	99	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.07
chr05	16562900	2+0-	chr05	16563068	1+3-	DEL	96	39	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	2.54
chr05	16570284	4+0-	chr05	16570300	4+0-	INV	-131	78	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	16698167	2+2-	chr05	16698392	1+3-	DEL	117	44	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	4.21
chr05	16787873	5+1-	chr05	16787933	5+1-	INV	-182	70	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	16829561	18+0-	chr05	16829835	0+18-	DEL	277	99	18	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|18	NA
chr05	16871480	0+2-	chr05	16872675	0+2-	INV	1018	73	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	1.04
chr05	16987325	8+0-	chr05	16987414	0+8-	DEL	98	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.74
chr05	17059769	15+0-	chr05	17060405	0+15-	DEL	633	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	0.02
chr05	14365254	4+1-	chr05	17465449	4+1-	INV	3099997	84	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	1.79
chr05	17163197	2+0-	chr05	17163327	0+2-	DEL	81	43	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	2.67
chr05	17205934	19+0-	chr05	17206894	0+19-	DEL	940	99	19	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|19	NA
chr05	17248456	10+0-	chr05	17248609	0+10-	DEL	141	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	0.32
chr05	17285723	7+0-	chr05	17286986	0+7-	DEL	1270	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	NA
chr05	17308342	2+0-	chr05	17308521	0+2-	DEL	87	60	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.35
chr05	17324762	6+0-	chr05	17325063	0+6-	DEL	220	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	NA
chr05	17333561	4+2-	chr05	17334366	0+4-	DEL	784	79	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.04
chr05	17456854	17+0-	chr05	17456998	0+17-	DEL	120	99	17	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|17	0.17
chr05	17473119	4+0-	chr05	17476303	0+4-	DEL	3122	86	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.01
chr05	17482594	17+0-	chr05	17482757	3+19-	DEL	134	99	16	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|16	0.46
chr05	17518558	7+0-	chr05	17519669	0+7-	DEL	1041	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	NA
chr05	17526913	14+0-	chr05	17527161	1+15-	DEL	247	99	14	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|14	NA
chr05	17529632	7+0-	chr05	17529927	0+7-	DEL	286	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	0.05
chr05	17579723	2+0-	chr05	17579833	0+2-	DEL	85	39	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	1.15
chr05	17646898	17+2-	chr05	17647836	12+14-	DEL	1087	99	14	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|14	1.19
chr05	17666462	14+0-	chr05	17667513	0+14-	DEL	1063	99	14	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|14	NA
chr05	17681323	15+0-	chr05	17682301	0+15-	DEL	952	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	0.07
chr05	17712728	19+1-	chr05	17713190	0+19-	DEL	507	99	19	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|19	0.03
chr05	17724591	3+0-	chr05	17726421	0+2-	DEL	1739	42	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	17727411	15+0-	chr05	17737895	0+15-	DEL	10438	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	0.00
chr05	17780188	6+0-	chr05	17780405	0+6-	DEL	181	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.24
chr05	17785970	12+0-	chr05	17795389	0+13-	DEL	9385	99	12	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|12	NA
chr05	17802206	4+0-	chr05	17802665	0+4-	DEL	386	88	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	NA
chr05	17843273	4+0-	chr05	17843605	0+2-	DEL	241	52	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.08
chr05	17846469	6+0-	chr05	17848345	0+6-	DEL	1865	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	3.79
chr05	17917967	7+0-	chr05	17918223	0+7-	DEL	243	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	0.21
chr05	17918753	18+0-	chr05	17919021	0+18-	DEL	260	99	18	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|18	0.10
chr05	17935193	2+0-	chr05	17935382	0+3-	DEL	87	54	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	2.17
chr05	17941409	3+0-	chr05	17941594	0+3-	DEL	109	74	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	4.97
chr05	17958270	1+2-	chr05	17959084	1+3-	INV	624	64	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	1.50
chr05	17994437	9+0-	chr05	17994882	0+9-	DEL	396	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	0.19
chr05	18026812	9+0-	chr05	18027031	0+9-	DEL	204	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	0.18
chr05	18034125	2+2-	chr05	18034397	4+2-	INV	51	72	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	4.50
chr05	18038427	0+4-	chr05	18038505	0+4-	INV	-80	68	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	18193652	6+0-	chr05	18193919	0+6-	DEL	201	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.30
chr05	18278717	14+0-	chr05	18290280	0+14-	DEL	11548	99	14	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|14	0.01
chr05	18298102	12+1-	chr05	18302014	0+12-	DEL	3894	99	12	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|12	0.04
chr05	18305776	3+0-	chr05	18306813	0+3-	DEL	1018	55	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.03
chr05	18327840	20+1-	chr05	18332246	0+19-	DEL	4405	99	19	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|19	0.01
chr05	18385694	2+0-	chr05	18395226	0+2-	DEL	9436	62	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	18407979	6+0-	chr05	18408292	0+6-	DEL	231	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	NA
chr05	18442569	17+0-	chr05	18443144	2+19-	DEL	585	99	17	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|17	0.02
chr05	18455033	21+0-	chr05	18455295	0+21-	DEL	254	99	21	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|21	NA
chr05	18569715	2+0-	chr05	18569881	0+2-	DEL	84	54	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	1.66
chr05	18572171	7+0-	chr05	18572557	0+7-	DEL	373	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	0.18
chr05	18596281	8+0-	chr05	18607084	0+10-	DEL	10775	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.00
chr05	18693046	1+4-	chr05	18693100	1+4-	INV	-93	71	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	18699495	2+0-	chr05	18700869	1+2-	DEL	1284	45	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.04
chr05	18742305	2+2-	chr05	18742501	1+1-	INV	78	57	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	1.38
chr05	18746143	17+0-	chr05	18746400	0+17-	DEL	265	99	17	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|17	NA
chr05	18747487	13+0-	chr05	18747939	1+14-	DEL	449	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	NA
chr05	18770973	6+2-	chr05	18771402	5+0-	INV	452	99	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	2.36
chr05	18803301	7+0-	chr05	18803554	0+7-	DEL	215	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	0.16
chr05	18831288	2+0-	chr05	18831452	0+2-	DEL	88	51	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	1.07
chr05	18855088	21+0-	chr05	18859492	0+20-	DEL	4418	99	20	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|20	NA
chr05	18936345	18+0-	chr05	18936602	0+18-	DEL	252	99	18	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|18	NA
chr05	18943560	3+0-	chr05	18944698	0+3-	DEL	1056	75	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.01
chr05	18994663	4+4-	chr05	18994987	4+4-	DEL	88	57	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	NA
chr05	19026401	4+0-	chr05	19026457	4+0-	INV	-91	71	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	19027130	7+0-	chr05	19027185	7+0-	INV	-98	98	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	NA
chr05	19028789	4+0-	chr05	19028883	0+4-	DEL	83	69	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	2.24
chr05	19172213	6+0-	chr05	19177530	0+6-	DEL	5312	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.00
chr05	19261419	2+0-	chr05	19261555	0+2-	DEL	97	41	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	5.15
chr05	19264651	4+0-	chr05	19264817	1+3-	DEL	80	41	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	1.21
chr05	19271231	7+0-	chr05	19271387	0+7-	DEL	102	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	1.19
chr05	19327746	4+1-	chr05	19327891	0+4-	DEL	89	75	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.84
chr05	19328571	9+0-	chr05	19329066	0+9-	DEL	443	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	0.11
chr05	19385480	18+0-	chr05	19385615	0+18-	DEL	132	99	18	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|18	0.27
chr05	19407494	3+0-	chr05	19407734	2+4-	DEL	317	53	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	NA
chr05	19408520	2+0-	chr05	19409235	0+2-	DEL	645	49	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	19660273	2+0-	chr05	19660737	10+12-	DEL	363	31	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.12
chr05	19416080	14+0-	chr05	19416221	0+14-	DEL	140	99	14	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|14	0.09
chr05	19418161	11+0-	chr05	19422626	0+11-	DEL	4449	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	NA
chr05	19447807	10+0-	chr05	19448762	1+10-	DEL	967	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	0.02
chr05	19463894	2+0-	chr05	19464043	0+2-	DEL	86	47	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	1.90
chr05	19476364	7+0-	chr05	19477080	0+7-	DEL	707	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	NA
chr05	19494053	10+0-	chr05	19494275	1+10-	DEL	209	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	0.06
chr05	19594832	3+0-	chr05	19606514	1+3-	DEL	11719	50	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	NA
chr05	19608947	8+0-	chr05	19609076	0+8-	DEL	122	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.46
chr05	19625679	6+0-	chr05	19627335	0+6-	DEL	1598	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.02
chr05	19628598	10+0-	chr05	19628780	0+10-	DEL	120	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	0.35
chr05	19647330	3+0-	chr05	19648022	0+3-	DEL	610	77	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.31
chr05	19655876	17+0-	chr05	19656227	0+17-	DEL	350	99	16	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|16	NA
chr05	19694476	4+2-	chr05	19694577	4+2-	INV	-85	66	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	19734086	13+0-	chr05	19734232	0+13-	DEL	103	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	0.34
chr05	19776046	16+0-	chr05	19776180	0+16-	DEL	110	99	16	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|16	0.36
chr05	19779396	4+1-	chr05	19779521	0+4-	DEL	83	78	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	1.14
chr05	19846895	11+0-	chr05	19847238	0+11-	DEL	349	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	NA
chr05	19860704	19+0-	chr05	19867949	1+20-	DEL	7239	99	19	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|19	NA
chr05	19909468	4+0-	chr05	19915983	0+4-	DEL	6430	96	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.02
chr05	19916549	5+0-	chr05	19920033	0+5-	DEL	3435	97	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.03
chr05	19968020	9+0-	chr05	19968233	0+9-	DEL	218	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	0.06
chr05	19971983	4+0-	chr05	19972095	0+4-	DEL	88	73	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	2.48
chr05	20000289	6+0-	chr05	20000950	0+6-	DEL	635	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.04
chr05	20002481	12+0-	chr05	20003406	0+12-	DEL	911	99	12	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|12	0.05
chr05	20059710	11+0-	chr05	20072624	0+11-	DEL	12924	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	0.00
chr05	20132643	15+0-	chr05	20145359	0+15-	DEL	12716	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	NA
chr05	20163469	4+0-	chr05	20163495	4+0-	INV	-121	76	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	20214040	24+0-	chr05	20222419	0+24-	DEL	8390	99	24	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|24	NA
chr05	20301209	2+0-	chr05	20301334	0+2-	DEL	102	39	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.95
chr05	20371710	17+0-	chr05	20374476	0+17-	DEL	2772	99	17	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|17	NA
chr05	20375546	18+0-	chr05	20375815	0+18-	DEL	259	99	18	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|18	NA
chr05	20466547	13+1-	chr05	20466663	0+12-	DEL	123	99	12	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|12	0.10
chr05	20478132	12+0-	chr05	20479299	0+12-	DEL	1124	99	12	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|12	0.01
chr05	20522821	13+0-	chr05	20522935	0+13-	DEL	95	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	0.71
chr05	20528873	5+0-	chr05	20534461	0+5-	DEL	5520	99	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	NA
chr05	20583909	0+3-	chr05	20584709	2+2-	INV	320	99	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	1.56
chr05	20608867	15+0-	chr05	20609131	0+15-	DEL	238	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	0.15
chr05	20640941	21+1-	chr05	20644342	0+20-	DEL	3413	99	20	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|20	NA
chr05	20681473	7+1-	chr05	20681528	7+1-	INV	-93	98	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	NA
chr05	20682142	3+0-	chr05	20682330	3+8-	DEL	101	56	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	2.32
chr05	20718086	6+0-	chr05	20718190	0+7-	DEL	89	98	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	1.09
chr05	20727808	11+0-	chr05	20728070	0+11-	DEL	242	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	0.15
chr05	20772847	4+4-	chr05	20772962	4+4-	INV	-59	65	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	20788403	22+0-	chr05	20788704	0+22-	DEL	300	99	22	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|22	NA
chr05	20922099	5+0-	chr05	20922553	0+5-	DEL	367	99	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.06
chr05	21001477	17+0-	chr05	21001635	0+17-	DEL	140	99	17	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|17	0.16
chr05	21005525	4+1-	chr05	21005692	4+1-	INV	-16	97	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	2.03
chr05	21019212	11+0-	chr05	21031618	0+13-	DEL	12399	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	0.00
chr05	21075008	30+0-	chr05	21075238	0+30-	DEL	232	99	30	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|30	0.11
chr05	21113867	5+9-	chr05	21113938	1+5-	DEL	217	58	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	2.29
chr05	21145948	3+0-	chr05	21146610	0+3-	DEL	598	66	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.11
chr05	21151909	2+0-	chr05	21157083	0+4-	DEL	5091	41	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.41
chr05	21218458	14+0-	chr05	21222143	0+14-	DEL	3689	99	14	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|14	0.00
chr05	21260549	11+1-	chr05	21262426	0+10-	DEL	1850	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	0.02
chr05	21280632	30+2-	chr05	21291708	1+29-	DEL	11085	99	28	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|28	NA
chr05	21431873	4+1-	chr05	21432012	0+3-	DEL	90	60	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.52
chr05	21437437	5+2-	chr05	21450180	0+5-	DEL	12684	84	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.00
chr05	21458066	6+0-	chr05	21458205	0+6-	DEL	98	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.61
chr05	21531482	14+0-	chr05	21548585	0+14-	DEL	17070	99	14	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|14	0.00
chr05	21554021	12+2-	chr05	21554403	0+11-	DEL	368	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	NA
chr05	21605888	16+0-	chr05	21606254	0+16-	DEL	370	99	16	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|16	NA
chr05	21613995	11+0-	chr05	21615166	0+11-	DEL	1138	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	0.03
chr05	21619766	6+0-	chr05	21619849	0+6-	DEL	93	98	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.64
chr05	21313025	4+0-	chr05	22034305	0+3-	DEL	721266	59	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	1.98
chr05	21763634	11+0-	chr05	21763873	0+11-	DEL	205	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	0.50
chr05	21772095	5+0-	chr05	21779347	0+5-	DEL	7170	99	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.02
chr05	21804902	10+0-	chr05	21817875	0+9-	DEL	12918	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	0.00
chr05	21829352	11+0-	chr05	21829617	0+11-	DEL	256	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	0.10
chr05	21862703	3+0-	chr05	21872881	0+3-	DEL	10109	70	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.01
chr05	21902682	3+0-	chr05	21902796	0+3-	DEL	87	55	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.61
chr05	21911758	2+0-	chr05	21911928	0+2-	DEL	85	56	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	1.19
chr05	21930273	0+6-	chr05	21930324	0+6-	INV	-96	99	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	NA
chr05	21941572	6+0-	chr05	21941868	0+6-	DEL	252	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	NA
chr05	22035003	3+0-	chr05	22035160	0+3-	DEL	86	70	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	3.32
chr05	22110265	8+0-	chr05	22110375	0+8-	DEL	99	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.94
chr05	22124939	4+0-	chr05	22125100	0+4-	DEL	115	77	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.39
chr05	22167180	12+0-	chr05	22173845	0+12-	DEL	6650	99	12	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|12	0.05
chr05	22235591	7+0-	chr05	22236066	0+7-	DEL	394	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	NA
chr05	22283453	0+4-	chr05	22283496	0+4-	INV	-104	73	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	22337432	4+0-	chr05	22349962	1+4-	DEL	12523	63	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	NA
chr05	22366185	6+0-	chr05	22367187	1+5-	DEL	969	67	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.10
chr05	22390298	3+0-	chr05	22390467	3+0-	INV	-15	99	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	3.87
chr05	22415588	6+0-	chr05	22423472	0+6-	DEL	7816	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.00
chr05	22461718	19+0-	chr05	22462054	0+19-	DEL	323	99	19	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|19	0.04
chr05	22596724	4+0-	chr05	22596940	0+4-	DEL	192	67	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.06
chr05	22609519	14+0-	chr05	22615442	0+14-	DEL	5936	99	14	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|14	0.01
chr05	22622450	7+0-	chr05	22622594	0+7-	DEL	115	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	0.08
chr05	22685673	3+0-	chr05	22685920	2+2-	INV	-35	83	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	1.35
chr05	22769645	9+0-	chr05	22769738	0+9-	DEL	100	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	0.12
chr05	22848166	18+0-	chr05	22852219	0+16-	DEL	4051	99	16	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|16	NA
chr05	22982323	18+0-	chr05	22983273	0+18-	DEL	930	99	18	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|18	0.02
chr05	23043405	8+0-	chr05	23044133	0+8-	DEL	680	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.08
chr05	23146944	11+0-	chr05	23154622	0+11-	DEL	7666	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	NA
chr05	23167626	11+0-	chr05	23177121	0+11-	DEL	9479	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	0.00
chr05	23202835	14+0-	chr05	23203082	0+14-	DEL	247	99	14	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|14	0.11
chr05	23221515	4+0-	chr05	23222016	0+4-	DEL	455	77	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.31
chr05	23223226	6+0-	chr05	23229356	0+6-	DEL	6079	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	NA
chr05	23322659	8+0-	chr05	23322802	0+8-	DEL	138	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.09
chr05	23323764	13+0-	chr05	23338430	0+13-	DEL	14647	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	0.00
chr05	23367286	5+0-	chr05	23372477	4+5-	DEL	5192	84	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	NA
chr05	23389725	14+0-	chr05	23392934	0+14-	DEL	3194	99	14	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|14	0.01
chr05	23423792	0+4-	chr05	23423855	0+4-	INV	-84	70	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	23437197	17+0-	chr05	23437875	0+17-	DEL	637	99	17	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|17	NA
chr05	23514546	6+0-	chr05	23514737	1+6-	DEL	244	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.20
chr05	23551792	15+0-	chr05	23556200	0+15-	DEL	4405	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	0.00
chr05	23563858	3+0-	chr05	23571705	0+3-	DEL	7780	68	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.04
chr05	23654949	2+1-	chr05	23655226	1+2-	DEL	169	57	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	4.53
chr05	23698371	15+0-	chr05	23698564	0+15-	DEL	166	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	0.27
chr05	23879033	2+0-	chr05	23879147	0+2-	DEL	80	41	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	1.22
chr05	23887788	8+0-	chr05	23889005	0+9-	DEL	1156	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	NA
chr05	23912772	13+1-	chr05	23913023	0+12-	DEL	259	99	12	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|12	0.16
chr05	23960076	15+0-	chr05	23972694	0+15-	DEL	12618	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	0.00
chr05	23998147	11+0-	chr05	23998525	0+11-	DEL	368	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	0.07
chr05	24039778	11+2-	chr05	24040322	2+9-	DEL	516	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	0.50
chr05	24050385	3+0-	chr05	24055775	0+4-	DEL	5302	63	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	NA
chr05	24064408	0+5-	chr05	24064478	0+5-	INV	-77	69	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	444151	2+1-	chr05	24315231	1+3-	DEL	23871058	47	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	1.98
chr05	24187912	6+0-	chr05	24188548	0+6-	DEL	552	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.09
chr05	24193947	6+0-	chr05	24194350	0+6-	DEL	334	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	NA
chr05	24221631	8+1-	chr05	24226111	0+8-	DEL	4468	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.01
chr05	24226944	10+0-	chr05	24227456	0+10-	DEL	476	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	0.06
chr05	24316521	7+1-	chr05	24316644	7+1-	INV	-24	89	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	NA
chr05	24326433	7+0-	chr05	24326540	0+7-	DEL	88	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	1.93
chr05	24346566	2+0-	chr05	24346727	0+2-	DEL	100	46	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	1.09
chr05	24362646	16+1-	chr05	24364914	0+16-	DEL	2255	99	16	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|16	0.01
chr05	24370172	11+0-	chr05	24370328	0+11-	DEL	123	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	0.16
chr05	24434788	15+0-	chr05	24440248	0+15-	DEL	5459	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	0.01
chr05	24647199	39+32-	chr05	24647923	27+38-	DEL	1047	99	38	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|38	0.90
chr05	24459922	13+0-	chr05	24460609	0+12-	DEL	674	99	12	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|12	NA
chr05	24461646	5+0-	chr05	24461728	0+5-	DEL	92	83	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.65
chr05	24572597	4+0-	chr05	24576808	0+4-	DEL	4119	99	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.03
chr05	24586683	3+0-	chr05	24587039	0+3-	DEL	350	52	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.04
chr05	24610822	9+0-	chr05	24610918	1+10-	DEL	92	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	0.23
chr05	24636977	1+2-	chr05	24637139	0+2-	INV	25	65	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.08
chr05	24657781	3+0-	chr05	24661751	0+3-	DEL	3935	56	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.01
chr05	24694331	4+0-	chr05	24694525	3+0-	INV	37	84	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	2.39
chr05	24720347	3+0-	chr05	24720556	0+3-	DEL	116	88	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.93
chr05	24789672	4+1-	chr05	24789759	0+4-	DEL	95	66	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.25
chr05	24807301	17+0-	chr05	24813032	1+16-	DEL	5724	99	16	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|16	0.01
chr05	24858291	6+3-	chr05	24858497	0+4-	DEL	138	85	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	NA
chr05	24871765	16+1-	chr05	24872748	1+16-	DEL	967	99	16	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|16	0.04
chr05	24914810	14+0-	chr05	24924035	0+14-	DEL	9202	99	14	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|14	0.15
chr05	24928722	3+0-	chr05	24953050	16+3-	DEL	24276	51	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.01
chr05	24968582	10+1-	chr05	24968955	0+9-	DEL	287	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	0.26
chr05	24975017	8+0-	chr05	24986355	0+8-	DEL	11307	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.00
chr05	25016149	6+0-	chr05	25016251	0+6-	DEL	92	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	1.88
chr05	25045702	4+0-	chr05	25052451	5+4-	DEL	6749	75	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.01
chr05	25149632	3+1-	chr05	25149822	0+2-	DEL	92	51	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	3.98
chr05	25165281	8+2-	chr05	25165406	0+6-	DEL	98	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.19
chr05	25197355	17+0-	chr05	25201913	0+17-	DEL	4542	99	17	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|17	0.01
chr05	25238098	14+1-	chr05	25251095	0+12-	DEL	13020	99	12	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|12	NA
chr05	25366909	21+2-	chr05	25378792	2+22-	DEL	11961	99	21	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|21	0.25
chr05	25405116	14+0-	chr05	25405451	0+14-	DEL	327	99	14	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|14	NA
chr05	25416530	19+0-	chr05	25429232	0+19-	DEL	12703	99	19	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|19	0.00
chr05	25434049	5+0-	chr05	25435444	0+5-	DEL	1297	99	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.01
chr05	25438728	2+2-	chr05	25438878	2+2-	INV	-123	62	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	25458317	10+0-	chr05	25458515	2+11-	DEL	164	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	0.39
chr05	25511344	8+0-	chr05	25511449	1+8-	DEL	83	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	1.41
chr05	25535018	25+0-	chr05	25535273	0+25-	DEL	244	99	25	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|25	0.05
chr05	25535758	11+0-	chr05	25535887	0+11-	DEL	96	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	1.02
chr05	25591409	15+0-	chr05	25606055	0+15-	DEL	14647	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	0.00
chr05	25672152	11+0-	chr05	25672383	0+11-	DEL	219	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	0.11
chr05	25673580	4+0-	chr05	25673673	0+4-	DEL	92	65	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	1.66
chr05	25693864	3+0-	chr05	25694055	0+3-	DEL	100	79	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	1.21
chr05	25709071	1+7-	chr05	25709194	1+7-	INV	-25	89	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	NA
chr05	25759271	5+0-	chr05	25759562	0+5-	DEL	225	99	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.56
chr05	25759962	10+0-	chr05	25760281	0+10-	DEL	294	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	0.04
chr05	25839766	0+4-	chr05	25839770	0+4-	INV	-142	82	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	25842393	7+1-	chr05	25842759	3+10-	DEL	347	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	0.15
chr05	25859640	12+0-	chr05	25872742	0+12-	DEL	13061	99	12	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|12	NA
chr05	26191687	3+2-	chr05	26192053	6+3-	DEL	498	43	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	NA
chr05	25911112	5+0-	chr05	25911303	0+5-	DEL	126	99	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.20
chr05	25957381	8+0-	chr05	25961009	0+8-	DEL	3574	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.04
chr05	25963764	13+0-	chr05	25964001	0+12-	DEL	227	99	12	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|12	0.11
chr05	25967441	4+0-	chr05	25967503	4+0-	INV	-85	70	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	25983756	25+0-	chr05	25996239	0+25-	DEL	12489	99	25	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|25	0.00
chr05	26014738	3+0-	chr05	26014877	0+3-	DEL	82	63	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.26
chr05	26018808	5+0-	chr05	26018886	0+5-	DEL	89	81	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.81
chr05	26032408	10+0-	chr05	26048065	0+10-	DEL	15657	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	0.01
chr05	26097361	22+0-	chr05	26097583	0+22-	DEL	209	99	22	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|22	NA
chr05	26098666	4+0-	chr05	26098693	4+0-	INV	-120	76	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	26148597	4+0-	chr05	26152027	0+4-	DEL	3381	78	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	NA
chr05	26187552	9+0-	chr05	26187629	0+9-	DEL	89	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	0.95
chr05	26203022	6+0-	chr05	26203231	3+5-	DEL	139	99	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.44
chr05	26206730	4+0-	chr05	26211609	0+5-	DEL	4828	77	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	2.07
chr05	26218124	10+0-	chr05	26223637	2+10-	DEL	5489	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	0.00
chr05	26229984	8+2-	chr05	26230937	0+6-	DEL	874	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	NA
chr05	26237413	0+5-	chr05	26237493	0+5-	INV	-125	68	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	26249244	16+0-	chr05	26249486	0+18-	DEL	247	99	16	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|16	NA
chr05	26264948	18+0-	chr05	26269511	0+18-	DEL	4545	99	18	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|18	0.01
chr05	26272675	10+0-	chr05	26272905	0+10-	DEL	216	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	NA
chr05	26283860	6+0-	chr05	26284391	0+6-	DEL	525	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.16
chr05	26321102	10+0-	chr05	26321257	0+10-	DEL	117	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	0.56
chr05	26352393	15+1-	chr05	26352746	1+15-	DEL	358	99	14	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|14	0.08
chr05	26353260	17+0-	chr05	26353633	0+15-	DEL	347	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	0.22
chr05	26363583	4+0-	chr05	26363702	0+4-	DEL	91	74	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	1.78
chr05	26411871	4+1-	chr05	26413023	0+4-	DEL	1084	90	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.01
chr05	26423550	19+0-	chr05	26434817	0+19-	DEL	11270	99	19	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|19	0.00
chr05	26436891	13+0-	chr05	26461596	0+13-	DEL	24669	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	NA
chr05	26515353	13+0-	chr05	26515560	0+13-	DEL	155	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	NA
chr05	26522105	4+0-	chr05	26535136	0+2-	DEL	12950	53	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.00
chr05	26594033	4+0-	chr05	26594078	4+0-	INV	-102	73	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	26603327	11+0-	chr05	26603545	1+11-	DEL	216	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	0.06
chr05	26668728	18+0-	chr05	26675215	0+18-	DEL	6499	99	18	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|18	0.00
chr05	26712551	0+4-	chr05	26712575	0+4-	INV	-123	77	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	26735823	6+0-	chr05	26736097	1+7-	DEL	253	97	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.15
chr05	26742715	5+0-	chr05	26742890	0+5-	DEL	146	95	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.07
chr05	26743186	11+0-	chr05	26743846	0+11-	DEL	613	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	0.02
chr05	26787529	18+2-	chr05	26788428	0+19-	DEL	878	99	18	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|18	0.13
chr05	7304825	0+10-	chr05	27181384	0+9-	INV	19876360	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	1.92
chr05	26876442	10+0-	chr05	26876547	1+12-	DEL	108	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	0.54
chr05	26924515	19+0-	chr05	26924662	0+19-	DEL	154	99	19	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|19	0.17
chr05	27049396	2+0-	chr05	27049499	0+2-	DEL	82	38	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	1.43
chr05	27106999	4+0-	chr05	27115159	0+4-	DEL	8127	73	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.00
chr05	27121414	2+0-	chr05	27121727	0+2-	DEL	252	46	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.13
chr05	27209914	11+0-	chr05	27210117	1+11-	DEL	232	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	0.06
chr05	27213807	4+0-	chr05	27213858	4+0-	INV	-96	72	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	27439978	2+1-	chr05	27440057	2+2-	DEL	88	36	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	1.60
chr05	27267436	11+0-	chr05	27284306	5+11-	DEL	16839	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	NA
chr05	27284397	5+11-	chr05	27284581	0+5-	DEL	118	99	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.07
chr05	27298555	14+0-	chr05	27299321	0+14-	DEL	749	99	14	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|14	0.04
chr05	27327409	11+2-	chr05	27330592	2+11-	DEL	3185	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	0.00
chr05	27331615	11+1-	chr05	27343597	6+16-	DEL	11975	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	0.00
chr05	27347109	18+0-	chr05	27353564	0+18-	DEL	6441	99	18	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|18	0.01
chr05	27398811	7+0-	chr05	27399940	0+7-	DEL	1106	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	0.01
chr05	27491722	12+0-	chr05	27492988	0+12-	DEL	1269	99	12	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|12	0.01
chr05	27496412	7+0-	chr05	27497065	0+7-	DEL	648	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	0.02
chr05	27537556	16+0-	chr05	27539368	0+16-	DEL	1801	99	16	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|16	0.01
chr05	27566045	17+0-	chr05	27577267	0+17-	DEL	11224	99	16	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|16	0.00
chr05	27726104	23+0-	chr05	27726453	0+21-	DEL	341	99	21	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|21	0.28
chr05	27637013	9+9-	chr05	27637340	9+9-	DEL	90	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	NA
chr05	27653708	17+1-	chr05	27655128	0+16-	DEL	1425	99	16	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|16	NA
chr05	27732583	6+0-	chr05	27733093	0+6-	DEL	508	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	1.42
chr05	27735499	1+5-	chr05	27735591	1+5-	INV	-95	67	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	27794940	5+0-	chr05	27795115	0+5-	DEL	91	99	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	1.01
chr05	27811017	3+0-	chr05	27821165	0+3-	DEL	10059	82	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.01
chr05	27824485	4+0-	chr05	27824581	0+4-	DEL	88	69	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	2.09
chr05	27831898	12+0-	chr05	27832121	0+12-	DEL	218	99	12	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|12	NA
chr05	27868372	13+0-	chr05	27868444	0+13-	DEL	89	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	1.14
chr05	27920659	4+2-	chr05	27920902	18+1-	INV	-32	61	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	1.97
chr05	27920902	18+1-	chr05	27927277	0+15-	DEL	6374	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	NA
chr05	27927817	13+1-	chr05	27928273	0+13-	DEL	450	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	0.22
chr05	27962295	11+0-	chr05	27963407	0+11-	DEL	1100	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	0.04
chr05	27968494	3+2-	chr05	27968623	3+2-	INV	-96	63	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	28018623	6+0-	chr05	28018678	6+0-	INV	-92	98	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	NA
chr05	28066881	15+0-	chr05	28067247	0+15-	DEL	365	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	0.04
chr05	28134123	14+0-	chr05	28134481	1+15-	DEL	361	99	14	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|14	0.15
chr05	28138668	3+0-	chr05	28139772	0+3-	DEL	1011	79	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.08
chr05	28326043	21+8-	chr05	28326630	13+20-	DEL	808	99	20	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|20	0.02
chr05	28217498	0+4-	chr05	28217527	0+4-	INV	-118	75	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	28308688	0+4-	chr05	28308719	0+4-	INV	-116	75	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	28336207	0+4-	chr05	28336269	0+4-	INV	-85	70	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	28356846	0+7-	chr05	28392350	0+7-	INV	35328	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	3.27
chr05	28358490	8+0-	chr05	28391113	7+0-	INV	32461	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	3.15
chr05	28359754	14+0-	chr05	28360393	0+16-	DEL	633	99	14	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|14	0.05
chr05	28379499	7+0-	chr05	28385137	7+0-	INV	5460	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	1.78
chr05	28404793	14+0-	chr05	28411314	0+14-	DEL	6501	99	14	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|14	0.01
chr05	28413963	5+0-	chr05	28415197	1+6-	DEL	1178	97	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.06
chr05	28417013	4+1-	chr05	28423485	0+3-	DEL	6432	60	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.01
chr05	28423989	6+1-	chr05	28424087	18+4-	DEL	98	56	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	1.03
chr05	28424249	18+4-	chr05	28440138	0+17-	DEL	15886	99	17	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|17	0.00
chr05	7136931	18+4-	chr05	28739087	0+18-	DEL	21602270	99	18	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|18	1.98
chr05	28570272	12+0-	chr05	28571109	0+12-	DEL	827	99	12	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|12	0.02
chr05	28571684	2+6-	chr05	28571976	2+6-	INV	-50	54	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	28661653	16+0-	chr05	28662691	0+16-	DEL	1004	99	16	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|16	0.08
chr05	28672239	4+0-	chr05	28673122	0+4-	DEL	839	80	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.02
chr05	28682127	25+0-	chr05	28682814	0+25-	DEL	697	99	25	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|25	0.02
chr05	28697720	9+0-	chr05	28697857	1+10-	DEL	215	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	NA
chr05	28706816	11+0-	chr05	28707868	0+11-	DEL	1029	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	0.03
chr05	28728840	2+0-	chr05	28728984	0+2-	DEL	91	44	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.76
chr05	28741110	10+0-	chr05	28741490	0+10-	DEL	373	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	0.04
chr05	28812411	23+0-	chr05	28812546	0+23-	DEL	139	99	23	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|23	0.09
chr05	28828267	0+4-	chr05	28828295	0+4-	INV	-154	86	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	28907763	4+0-	chr05	28907922	0+4-	DEL	95	84	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.70
chr05	28949340	8+1-	chr05	28949792	0+8-	DEL	523	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.03
chr05	28968212	4+1-	chr05	28968663	0+3-	DEL	357	68	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.06
chr05	29002504	3+0-	chr05	29002766	0+3-	DEL	178	71	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.20
chr05	29006964	11+0-	chr05	29010956	0+11-	DEL	3985	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	0.02
chr05	29042248	0+4-	chr05	29042382	0+4-	INV	-67	63	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	29050727	13+0-	chr05	29050902	0+13-	DEL	178	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	NA
chr05	29083087	4+0-	chr05	29092356	0+4-	DEL	9244	69	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	NA
chr05	29099686	10+0-	chr05	29099916	0+10-	DEL	195	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	0.23
chr05	29208370	11+1-	chr05	29208575	0+13-	DEL	172	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	NA
chr05	29216678	1+4-	chr05	29216822	1+4-	INV	-129	62	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	29275069	15+0-	chr05	29281508	0+14-	DEL	6455	99	14	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|14	0.00
chr05	29290599	4+0-	chr05	29290735	0+4-	DEL	85	82	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	1.15
chr05	29342588	24+1-	chr05	29343862	0+23-	DEL	1271	99	23	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|23	0.02
chr05	29348798	18+0-	chr05	29355187	3+19-	DEL	6425	99	18	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|18	NA
chr05	29379492	3+0-	chr05	29379594	0+3-	DEL	90	53	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	1.44
chr05	29390946	18+0-	chr05	29402051	1+18-	DEL	11110	99	18	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|18	NA
chr05	29406589	4+4-	chr05	29406917	4+4-	DEL	87	56	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	NA
chr05	29410339	16+2-	chr05	29411515	0+15-	DEL	1193	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	0.01
chr05	29427167	5+0-	chr05	29432415	1+11-	DEL	5163	99	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.04
chr05	29431819	0+6-	chr05	29432511	1+11-	INV	485	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.08
chr05	29446227	13+1-	chr05	29447628	0+12-	DEL	1378	99	12	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|12	NA
chr05	29450468	9+0-	chr05	29451503	0+10-	DEL	1022	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	0.03
chr05	29506556	3+1-	chr05	29506890	0+3-	DEL	247	60	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.16
chr05	29729809	4+0-	chr05	29729951	4+0-	INV	-43	62	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr05	29742845	0+2-	chr05	29743032	0+2-	INV	-2	75	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	2.67
chr10	63809	16+0-	chr10	63929	0+17-	DEL	110	99	16	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|16	0.49
chr10	93873	18+0-	chr10	94148	0+18-	DEL	266	99	18	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|18	0.10
chr10	172296	6+0-	chr10	172531	0+6-	DEL	165	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.23
chr10	174683	17+0-	chr10	174823	0+17-	DEL	112	99	17	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|17	0.09
chr10	179245	2+4-	chr10	179322	2+4-	INV	-154	68	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr10	288971	15+0-	chr10	289241	1+15-	DEL	252	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	0.25
chr10	316433	6+0-	chr10	316543	6+0-	INV	-77	65	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr10	316578	6+0-	chr10	318111	0+2-	DEL	1475	38	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.02
chr10	337453	9+0-	chr10	337698	0+9-	DEL	226	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	0.11
chr10	338171	3+0-	chr10	338647	0+3-	DEL	428	59	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	NA
chr10	346275	3+0-	chr10	346543	0+3-	DEL	188	75	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.20
chr10	447346	0+4-	chr10	447430	0+4-	INV	-77	67	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr10	577998	4+2-	chr10	579106	2+0-	INV	1124	57	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	3.48
chr10	577998	4+2-	chr10	579382	1+3-	INV	1329	58	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	4.21
chr10	583302	5+0-	chr10	583930	0+5-	DEL	597	87	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.02
chr10	660720	13+0-	chr10	664406	0+13-	DEL	3662	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	NA
chr10	731442	13+0-	chr10	731771	2+13-	DEL	342	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	NA
chr10	744791	8+0-	chr10	745136	1+8-	DEL	256	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	0.08
chr10	807020	13+1-	chr10	807617	0+12-	DEL	603	99	12	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|12	0.07
chr10	838987	14+0-	chr10	839168	0+14-	DEL	150	99	14	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|14	0.14
chr10	847612	0+4-	chr10	847801	0+4-	INV	-16	99	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.75
chr10	850967	6+0-	chr10	851680	0+6-	DEL	690	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	NA
chr10	954435	8+0-	chr10	955933	0+6-	DEL	1488	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.03
chr10	879697	10+0-	chr10	879963	0+10-	DEL	257	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	NA
chr10	909148	4+0-	chr10	909186	4+0-	INV	-109	74	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr10	935669	19+0-	chr10	935903	0+19-	DEL	220	99	19	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|19	0.06
chr10	1039708	10+0-	chr10	1047870	2+12-	DEL	8153	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	0.00
chr10	1050495	8+0-	chr10	1056369	0+8-	DEL	5832	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	NA
chr10	1081201	7+0-	chr10	1082269	0+7-	DEL	1013	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	NA
chr10	1120334	5+0-	chr10	1121634	0+5-	DEL	1290	85	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	NA
chr10	1143299	15+0-	chr10	1154603	1+16-	DEL	11311	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	NA
chr10	1185843	17+0-	chr10	1189426	0+17-	DEL	3585	99	17	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|17	0.01
chr10	1215971	13+0-	chr10	1222487	0+13-	DEL	6491	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	0.01
chr10	1245641	3+0-	chr10	1264793	1+4-	DEL	19056	88	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	NA
chr10	1266544	2+2-	chr10	1267134	0+2-	DEL	515	40	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.05
chr10	1383675	13+0-	chr10	1383773	0+13-	DEL	98	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	0.80
chr10	1407209	12+1-	chr10	1416992	0+11-	DEL	9801	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	NA
chr10	1472396	21+0-	chr10	1472892	0+21-	DEL	484	99	21	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|21	0.20
chr10	1477084	5+0-	chr10	1477485	0+5-	DEL	324	99	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.31
chr10	1481449	2+0-	chr10	1481632	0+2-	DEL	117	48	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	1.39
chr10	1482144	4+0-	chr10	1493136	1+4-	DEL	10980	70	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.00
chr10	1496254	10+0-	chr10	1496479	0+10-	DEL	161	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	0.53
chr10	1497015	9+0-	chr10	1498148	0+9-	DEL	1105	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	0.03
chr10	1536412	5+1-	chr10	1536602	0+5-	DEL	135	89	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.07
chr10	1536834	3+0-	chr10	1537108	1+3-	DEL	178	82	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.49
chr10	1548657	4+0-	chr10	1557434	0+4-	DEL	8694	96	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.01
chr10	1559823	4+0-	chr10	1560106	0+4-	DEL	222	82	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.05
chr10	1570992	4+0-	chr10	1574715	0+4-	DEL	3665	90	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.02
chr10	1583919	15+0-	chr10	1584888	0+15-	DEL	957	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	0.02
chr10	1602892	14+0-	chr10	1603115	2+16-	DEL	198	99	14	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|14	0.47
chr10	1621215	7+0-	chr10	1622037	0+7-	DEL	739	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	0.05
chr10	1674106	3+2-	chr10	1674553	0+5-	DEL	430	58	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	6.59
chr10	1707368	10+1-	chr10	1708749	0+10-	DEL	1357	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	0.05
chr10	1758141	11+0-	chr10	1762880	1+11-	DEL	4739	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	0.00
chr10	1772776	11+0-	chr10	1772863	0+11-	DEL	102	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	0.12
chr10	1787765	7+0-	chr10	1789262	3+7-	DEL	1461	63	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	2.72
chr10	1794384	13+8-	chr10	1794578	13+0-	INV	171	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	0.46
chr10	1794384	13+8-	chr10	1798689	0+9-	INV	4132	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.07
chr10	1805822	6+0-	chr10	1811617	0+9-	DEL	5730	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.00
chr10	1818199	5+0-	chr10	1819463	0+5-	DEL	1251	89	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.02
chr10	1879274	5+0-	chr10	1887602	0+5-	DEL	8256	99	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.00
chr10	2056980	4+0-	chr10	2057444	0+4-	DEL	467	67	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	NA
chr10	2067697	8+0-	chr10	2068034	0+8-	DEL	264	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.04
chr10	2085609	4+0-	chr10	2085824	0+3-	DEL	179	68	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.18
chr10	2087974	4+0-	chr10	2088248	0+4-	DEL	243	73	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.25
chr10	2102571	6+0-	chr10	2103095	0+6-	DEL	440	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.11
chr10	2109687	15+0-	chr10	2109998	0+15-	DEL	277	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	0.13
chr10	2119191	13+0-	chr10	2122598	0+13-	DEL	3392	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	0.02
chr10	2145932	18+0-	chr10	2146453	0+16-	DEL	495	99	16	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|16	NA
chr10	2152645	0+3-	chr10	2240933	0+3-	INV	88111	99	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	1.45
chr10	2154284	19+2-	chr10	2154642	0+19-	DEL	468	99	19	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|19	0.12
chr10	2189980	13+0-	chr10	2190638	0+13-	DEL	613	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	0.02
chr10	2242712	6+0-	chr10	2243068	0+6-	DEL	268	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.04
chr10	2244435	5+0-	chr10	2244571	0+3-	DEL	153	56	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.09
chr10	2254391	7+0-	chr10	2254671	0+8-	DEL	251	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	NA
chr10	2262690	4+0-	chr10	2263111	0+3-	DEL	342	66	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.20
chr10	2275447	8+2-	chr10	2276221	0+8-	DEL	697	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.02
chr10	2552731	9+5-	chr10	2552869	3+8-	DEL	106	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	2.46
chr10	2279545	5+0-	chr10	2280236	0+5-	DEL	611	99	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.06
chr10	2317057	9+0-	chr10	2317700	0+9-	DEL	575	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	0.02
chr10	2346956	6+0-	chr10	2349775	0+6-	DEL	2808	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.04
chr10	2460953	15+0-	chr10	2512834	15+0-	INV	51695	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	1.83
chr10	2474194	2+1-	chr10	2475030	0+2-	DEL	758	41	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr10	2560007	0+3-	chr10	2560314	0+2-	INV	112	63	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	1.82
chr10	2574219	0+4-	chr10	2574327	0+4-	INV	-68	65	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr10	2576787	9+0-	chr10	2580793	0+12-	DEL	4007	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	0.00
chr10	2584597	14+0-	chr10	2584747	0+14-	DEL	154	99	14	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|14	0.08
chr10	2593515	5+0-	chr10	2593931	0+5-	DEL	319	99	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.07
chr10	2596922	10+0-	chr10	2598247	8+11-	DEL	1332	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	NA
chr10	2598409	8+11-	chr10	2598528	2+9-	DEL	111	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	0.10
chr10	2611952	8+0-	chr10	2618736	0+8-	DEL	6751	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.00
chr10	2622482	17+1-	chr10	2622716	0+16-	DEL	213	99	16	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|16	0.28
chr10	2978157	6+2-	chr10	2981621	0+6-	DEL	3609	69	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.47
chr10	2676441	20+0-	chr10	2681824	0+20-	DEL	5373	99	20	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|20	0.01
chr10	2714620	10+2-	chr10	2715632	0+10-	DEL	1062	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	0.06
chr10	2777062	9+0-	chr10	2777382	0+9-	DEL	295	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	0.04
chr10	2789377	7+0-	chr10	2789797	0+7-	DEL	435	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	0.03
chr10	2790745	11+0-	chr10	2791038	0+11-	DEL	273	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	0.05
chr10	2797284	2+0-	chr10	2797453	0+2-	DEL	86	54	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	2.16
chr10	2799992	8+0-	chr10	2800257	0+8-	DEL	277	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.05
chr10	2865038	16+0-	chr10	2866385	0+16-	DEL	1357	99	16	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|16	0.04
chr10	2886884	6+0-	chr10	2887294	0+7-	DEL	373	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.10
chr10	2892708	5+0-	chr10	2893973	1+5-	DEL	1264	83	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	NA
chr10	2901153	6+0-	chr10	2901417	0+6-	DEL	252	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.05
chr10	2924740	17+0-	chr10	2924887	0+17-	DEL	153	99	17	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|17	0.08
chr10	2927558	10+2-	chr10	2927702	0+10-	DEL	148	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	0.08
chr10	2929214	5+0-	chr10	2929395	0+5-	DEL	91	99	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.98
chr10	2931475	22+0-	chr10	2931691	0+22-	DEL	212	99	22	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|22	0.24
chr10	2952627	4+0-	chr10	2956084	0+4-	DEL	3363	99	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	NA
chr10	2971237	13+1-	chr10	2974253	0+13-	DEL	3013	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	0.04
chr10	2998372	2+0-	chr10	2999014	0+2-	DEL	562	53	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.13
chr10	3019776	2+0-	chr10	3020050	2+6-	INV	-42	99	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.54
chr10	3023077	2+0-	chr10	3023170	1+3-	DEL	86	37	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.59
chr10	3029958	9+0-	chr10	3031375	0+9-	DEL	1356	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	NA
chr10	3035155	3+0-	chr10	3035333	0+3-	DEL	84	84	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.43
chr10	3036102	6+0-	chr10	3036381	0+6-	DEL	248	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.19
chr10	3036765	6+0-	chr10	3036875	0+6-	DEL	88	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.94
chr10	3037919	7+0-	chr10	3038253	0+7-	DEL	313	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	NA
chr10	3043344	5+0-	chr10	3043576	0+5-	DEL	186	99	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.06
chr10	3058543	4+0-	chr10	3058850	0+4-	DEL	228	94	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	1.73
chr10	3059231	27+2-	chr10	3060055	0+29-	DEL	810	99	27	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|27	0.74
chr10	3084713	7+0-	chr10	3084900	0+7-	DEL	100	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	1.23
chr10	3086149	14+0-	chr10	3086843	0+14-	DEL	689	99	14	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|14	0.06
chr10	3088182	13+0-	chr10	3088729	0+10-	DEL	505	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	0.31
chr10	3094209	9+0-	chr10	3094380	0+9-	DEL	129	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	0.07
chr10	3104620	2+0-	chr10	3104792	3+2-	DEL	119	33	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.07
chr10	3357135	15+0-	chr10	3393347	15+0-	INV	35999	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	1.17
chr10	3427516	17+0-	chr10	3427757	0+17-	DEL	240	99	17	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|17	NA
chr10	3446833	23+1-	chr10	3458106	0+23-	DEL	11276	99	23	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|23	0.00
chr10	3475638	4+0-	chr10	3475736	0+4-	DEL	89	68	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.80
chr10	3477058	13+2-	chr10	3477407	2+13-	DEL	335	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	4.55
chr10	3583464	11+4-	chr10	3587416	0+7-	DEL	3938	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	NA
chr10	3591012	2+0-	chr10	3591181	0+2-	DEL	79	58	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.37
chr10	3644527	0+2-	chr10	3644696	0+2-	INV	-21	72	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	2.68
chr10	3657068	4+0-	chr10	3657235	0+3-	DEL	110	72	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	1.73
chr10	3677463	10+0-	chr10	3677558	0+10-	DEL	101	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	0.12
chr10	3694099	16+0-	chr10	3694201	3+16-	DEL	102	99	16	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|16	1.55
chr10	3694384	3+16-	chr10	3695574	0+3-	DEL	1117	51	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.50
chr10	3700160	2+0-	chr10	3700329	0+2-	DEL	94	51	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.22
chr10	3780038	4+0-	chr10	3780216	0+4-	DEL	98	96	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.14
chr10	3788195	6+1-	chr10	3789455	0+6-	DEL	1229	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	NA
chr10	3790652	6+0-	chr10	3792101	3+6-	DEL	1417	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	2.83
chr10	3795924	8+0-	chr10	3798503	0+8-	DEL	2522	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.06
chr10	3805046	18+0-	chr10	3805164	0+18-	DEL	118	99	18	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|18	0.10
chr10	3815984	2+0-	chr10	3823324	0+2-	DEL	7299	42	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.00
chr10	3828571	4+1-	chr10	3828732	0+3-	DEL	86	72	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	2.17
chr10	3862625	0+4-	chr10	3862647	0+4-	INV	-125	77	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr10	3961924	8+0-	chr10	3965644	0+8-	DEL	3655	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	NA
chr10	3970185	8+1-	chr10	3970375	7+7-	DEL	165	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	0.20
chr10	3970487	7+7-	chr10	3971037	0+7-	DEL	498	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	0.42
chr10	3972354	10+0-	chr10	3973368	0+10-	DEL	983	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	0.03
chr10	4038084	8+0-	chr10	4043212	0+8-	DEL	5104	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.00
chr10	4063384	10+0-	chr10	4074494	0+10-	DEL	11109	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	0.00
chr10	4081945	11+0-	chr10	4082443	0+11-	DEL	471	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	NA
chr10	4233360	5+0-	chr10	4233469	0+5-	DEL	88	90	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.11
chr10	4247082	2+0-	chr10	4248374	1+2-	DEL	1225	48	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr10	4249057	20+1-	chr10	4251079	0+19-	DEL	1997	99	19	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|19	0.01
chr10	4268080	3+0-	chr10	4271282	0+3-	DEL	3168	58	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.01
chr10	4300069	9+0-	chr10	4311143	0+9-	DEL	11079	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	NA
chr10	4320355	10+0-	chr10	4320850	0+10-	DEL	444	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	0.09
chr10	4327968	6+0-	chr10	4328196	0+6-	DEL	167	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.17
chr10	4385473	4+0-	chr10	4392454	0+4-	DEL	6936	77	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.01
chr10	4403836	8+0-	chr10	4404342	0+8-	DEL	481	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.11
chr10	4409924	10+0-	chr10	4410048	0+11-	DEL	97	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	0.86
chr10	4416173	20+0-	chr10	4417077	0+20-	DEL	910	99	20	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|20	0.03
chr10	4455844	15+0-	chr10	4466310	2+17-	DEL	10476	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	NA
chr10	4470120	22+0-	chr10	4473035	1+23-	DEL	2914	99	22	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|22	NA
chr10	4483092	17+0-	chr10	4488532	0+17-	DEL	5422	99	17	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|17	0.01
chr10	4521747	14+1-	chr10	4521816	0+13-	DEL	95	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	0.88
chr10	4849200	13+0-	chr10	4854325	8+13-	DEL	5137	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	0.01
chr10	4702540	8+0-	chr10	4703206	1+9-	DEL	643	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.04
chr10	4713948	19+0-	chr10	4725359	0+19-	DEL	11421	99	19	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|19	0.00
chr10	4763875	8+0-	chr10	4775586	0+10-	DEL	11681	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.00
chr10	4866162	11+0-	chr10	4866505	0+11-	DEL	341	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	NA
chr10	4887673	4+1-	chr10	4890740	0+4-	DEL	3064	70	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	NA
chr10	4899052	2+0-	chr10	4910765	0+2-	DEL	11683	40	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.02
chr10	4955424	3+0-	chr10	4961568	0+3-	DEL	6063	73	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	NA
chr10	5185652	5+0-	chr10	5188519	0+5-	DEL	2864	83	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.01
chr10	5190052	12+0-	chr10	5196373	0+12-	DEL	6305	99	12	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|12	0.01
chr10	5218132	3+0-	chr10	5219384	1+3-	DEL	1282	50	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.11
chr10	5356785	15+4-	chr10	5357229	0+15-	DEL	500	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	NA
chr10	5282280	19+0-	chr10	5283221	0+21-	DEL	918	99	19	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|19	0.03
chr10	5293216	5+0-	chr10	5293333	0+5-	DEL	90	92	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	1.10
chr10	5348122	7+0-	chr10	5355980	1+8-	DEL	7839	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	0.02
chr10	5360273	7+0-	chr10	5365249	0+7-	DEL	4955	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	0.26
chr10	5392629	5+1-	chr10	5412445	0+4-	DEL	19765	71	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.01
chr10	5417550	4+1-	chr10	5427207	0+4-	DEL	9678	68	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.06
chr10	5454584	3+0-	chr10	5457282	0+3-	DEL	2630	69	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	NA
chr10	5460690	17+9-	chr10	5460852	0+8-	DEL	104	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.15
chr10	5476672	8+0-	chr10	5483289	0+8-	DEL	6619	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	NA
chr10	5672401	4+0-	chr10	5675930	5+2-	INV	3346	85	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	3.63
chr10	5806092	10+2-	chr10	5806186	0+10-	DEL	94	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	0.24
chr10	5848151	2+0-	chr10	5860215	0+2-	DEL	12018	43	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.00
chr10	5921083	3+0-	chr10	5923734	0+6-	DEL	2572	60	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	NA
chr10	5950444	3+0-	chr10	5961784	0+3-	DEL	11287	58	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	NA
chr10	5969253	0+4-	chr10	5969293	0+4-	INV	-108	73	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr10	5969842	3+0-	chr10	6005830	0+2-	DEL	35954	45	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.00
chr10	6080065	19+0-	chr10	6080361	0+19-	DEL	298	99	19	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|19	0.05
chr10	6094287	9+1-	chr10	6094413	0+8-	DEL	88	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.75
chr10	6135342	8+0-	chr10	6136618	0+8-	DEL	1245	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.02
chr10	6152134	2+0-	chr10	6155668	0+2-	DEL	3459	51	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.03
chr10	6178026	13+0-	chr10	6186583	0+13-	DEL	8551	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	NA
chr10	6217483	13+0-	chr10	6232377	0+13-	DEL	14895	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	0.00
chr10	6259616	16+0-	chr10	6259804	0+16-	DEL	166	99	16	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|16	NA
chr10	6391605	12+0-	chr10	6402925	0+12-	DEL	11269	99	12	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|12	0.01
chr10	6408557	12+0-	chr10	6421466	3+13-	DEL	12965	99	12	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|12	0.00
chr10	6435864	11+0-	chr10	6447955	0+11-	DEL	12075	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	0.01
chr10	6548194	8+0-	chr10	6548652	0+8-	DEL	398	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.25
chr10	6638978	6+0-	chr10	6639223	0+6-	DEL	244	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.16
chr10	6647346	2+0-	chr10	6647565	0+2-	DEL	171	43	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.24
chr10	6693425	6+0-	chr10	6695536	0+6-	DEL	2069	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	NA
chr10	6703173	17+0-	chr10	6708360	0+17-	DEL	5161	99	17	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|17	0.03
chr10	6760760	4+0-	chr10	6760893	0+4-	DEL	87	78	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.63
chr10	6801603	17+0-	chr10	6812933	16+17-	DEL	11329	99	17	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|17	NA
chr10	6813177	16+17-	chr10	6836392	0+16-	DEL	23202	99	16	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|16	0.00
chr10	7305457	27+1-	chr10	7305626	6+27-	DEL	310	99	27	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|27	NA
chr10	6909419	2+2-	chr10	6909465	2+2-	INV	-141	72	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr10	6921752	3+0-	chr10	6924541	0+3-	DEL	2729	64	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	NA
chr10	6959377	4+0-	chr10	6974464	0+4-	DEL	15071	73	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.01
chr10	7020518	6+0-	chr10	7021167	5+0-	INV	454	99	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	3.09
chr10	7020706	0+11-	chr10	7021415	1+11-	INV	482	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	2.86
chr10	7113470	17+0-	chr10	7113837	0+17-	DEL	338	99	17	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|17	0.23
chr10	7141517	7+0-	chr10	7153042	0+7-	DEL	11516	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	0.00
chr10	7153953	2+0-	chr10	7217366	0+2-	DEL	63329	55	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.00
chr10	7222539	15+0-	chr10	7222666	0+15-	DEL	93	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	1.13
chr10	7228408	9+0-	chr10	7239761	0+11-	DEL	11317	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	0.00
chr10	7241095	7+0-	chr10	7241482	0+7-	DEL	353	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	3.78
chr10	7293017	9+0-	chr10	7293294	0+9-	DEL	277	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	NA
chr10	7316895	8+0-	chr10	7328882	0+8-	DEL	11962	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.01
chr10	7363571	19+0-	chr10	7369496	0+19-	DEL	5923	99	19	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|19	0.01
chr10	7397294	2+1-	chr10	7397667	4+2-	INV	55	76	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.60
chr10	578159	0+3-	chr10	7463348	0+4-	INV	6884937	70	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	1.33
chr10	7414347	2+0-	chr10	7414497	0+2-	DEL	86	47	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	2.13
chr10	7436502	10+1-	chr10	7437096	0+10-	DEL	525	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	0.05
chr10	7450095	14+0-	chr10	7450469	1+15-	DEL	346	99	14	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|14	0.11
chr10	7488379	6+0-	chr10	7494374	0+6-	DEL	5987	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.01
chr10	7560735	2+0-	chr10	7560905	0+2-	DEL	82	57	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	3.04
chr10	7582568	3+0-	chr10	7585099	0+3-	DEL	2491	59	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	NA
chr10	7600461	19+0-	chr10	7611765	0+19-	DEL	11309	99	19	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|19	NA
chr10	7613002	18+9-	chr10	7675888	18+9-	INV	62650	99	27	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|27	1.38
chr10	7659123	11+0-	chr10	7659278	0+10-	DEL	112	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	0.56
chr10	7695314	1+5-	chr10	7695470	1+5-	INV	-92	61	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr10	7702752	4+0-	chr10	7704284	0+4-	DEL	1535	64	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.01
chr10	7711388	14+1-	chr10	7715396	0+14-	DEL	3990	99	14	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|14	8.19
chr10	7712942	4+2-	chr10	7713109	4+2-	INV	-62	61	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr10	7801857	9+0-	chr10	7802585	0+9-	DEL	715	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	0.06
chr10	7809457	8+0-	chr10	7810136	0+8-	DEL	626	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.19
chr10	7815037	0+4-	chr10	7815088	0+4-	INV	-96	72	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr10	7965913	10+0-	chr10	7966476	1+10-	DEL	562	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	1.24
chr10	7984087	8+0-	chr10	7984711	0+8-	DEL	557	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.14
chr10	8038155	9+1-	chr10	8038988	0+8-	DEL	810	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	1.54
chr10	8039921	5+1-	chr10	8040256	0+5-	DEL	247	99	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.16
chr10	8288628	2+0-	chr10	8289001	0+2-	DEL	314	46	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.04
chr10	8293416	9+0-	chr10	8293676	1+9-	DEL	242	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	0.05
chr10	8296901	2+0-	chr10	8297220	0+2-	DEL	235	55	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.30
chr10	8371647	3+0-	chr10	8374885	0+3-	DEL	3163	69	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.00
chr10	8411418	4+0-	chr10	8416769	0+3-	DEL	5253	79	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.00
chr10	8430003	3+0-	chr10	8430184	0+3-	DEL	84	91	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.21
chr10	8431405	2+0-	chr10	8431607	2+2-	DEL	108	65	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	1.28
chr10	8431654	2+2-	chr10	8444145	0+4-	DEL	12452	49	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.00
chr10	8479463	8+0-	chr10	8490263	0+8-	DEL	10778	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.01
chr02	32853140	3+1-	chr10	8913625	3+8-	INV	-182	62	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	-19.09
chr10	8912686	4+1-	chr10	8913420	3+8-	DEL	705	57	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.04
chr10	8566113	5+0-	chr10	8569687	0+5-	DEL	3586	82	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	NA
chr10	8577404	10+1-	chr10	8585387	0+10-	DEL	7964	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	0.00
chr10	8598493	10+0-	chr10	8598855	0+10-	DEL	341	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	0.15
chr10	8643519	3+0-	chr10	8654327	0+3-	DEL	10717	82	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	NA
chr10	8664077	24+0-	chr10	8678579	0+23-	DEL	14509	99	23	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|23	0.00
chr10	8722365	4+0-	chr10	8759126	0+4-	DEL	36702	87	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	NA
chr10	8848856	5+0-	chr10	8867053	1+5-	DEL	18177	92	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	NA
chr10	8876789	10+0-	chr10	8886455	0+10-	DEL	9631	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	0.01
chr10	8966856	0+4-	chr10	8966865	0+4-	INV	-138	80	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr10	8970067	6+1-	chr10	8973483	0+6-	DEL	3399	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	NA
chr10	9043152	9+2-	chr10	9053926	1+10-	DEL	10807	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	0.00
chr10	9070653	4+9-	chr10	9072865	4+0-	INV	2201	99	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	3.10
chr10	9070653	4+9-	chr10	9073181	0+9-	INV	2346	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	2.74
chr10	9165024	3+0-	chr10	9165171	0+3-	DEL	83	66	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	2.17
chr10	9218506	20+0-	chr10	9226449	0+20-	DEL	7961	99	20	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|20	NA
chr10	9286374	17+2-	chr10	9288710	1+17-	DEL	2454	99	17	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|17	3.83
chr10	9291458	5+0-	chr10	9304383	1+6-	DEL	12921	78	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	NA
chr10	9314563	8+1-	chr10	9314925	0+7-	DEL	294	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	0.34
chr10	9394243	4+0-	chr10	9400639	0+4-	DEL	6299	99	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	1.34
chr10	9477260	4+0-	chr10	9490626	0+4-	DEL	13320	76	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.00
chr10	9504068	4+0-	chr10	9504224	0+4-	DEL	86	90	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.40
chr10	9543334	8+0-	chr10	9551039	9+8-	DEL	7692	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.01
chr10	9551277	9+8-	chr10	9551399	0+9-	DEL	103	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	0.19
chr10	9558445	9+0-	chr10	9558575	0+9-	DEL	95	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	0.64
chr10	9559402	4+0-	chr10	9559578	0+4-	DEL	83	99	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.94
chr10	9565596	0+4-	chr10	9565663	0+4-	INV	-80	69	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr10	9602670	11+0-	chr10	9603727	0+11-	DEL	1051	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	0.01
chr10	9630965	13+0-	chr10	9632446	0+13-	DEL	1453	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	0.11
chr10	9670510	15+0-	chr10	9671954	0+13-	DEL	1457	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	NA
chr10	9708990	19+0-	chr10	9712656	0+19-	DEL	3670	99	19	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|19	1.58
chr10	9713572	7+0-	chr10	9719651	0+7-	DEL	6063	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	0.01
chr10	9731963	3+0-	chr10	9743482	0+3-	DEL	11431	80	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.01
chr10	9784524	0+4-	chr10	9784589	0+4-	INV	-83	70	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr10	9804846	20+4-	chr10	9814106	0+20-	DEL	9259	99	20	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|20	NA
chr10	9815442	10+0-	chr10	9815769	0+10-	DEL	285	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	NA
chr10	9877327	5+1-	chr10	9891991	0+3-	DEL	14576	67	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.01
chr10	9911522	6+0-	chr10	9911641	0+6-	DEL	94	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.59
chr10	9924454	4+0-	chr10	9924508	4+0-	INV	-137	71	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr10	9947222	3+0-	chr10	9947353	0+3-	DEL	84	60	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	2.10
chr10	9800929	7+0-	chr10	10312289	0+7-	DEL	511295	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	1.50
chr10	10008070	13+0-	chr10	10008189	0+13-	DEL	103	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	0.39
chr10	10019266	3+0-	chr10	10029607	0+2-	DEL	10243	67	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr10	10075403	9+0-	chr10	10079029	0+9-	DEL	3589	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	0.01
chr10	10187153	2+0-	chr10	10187347	0+2-	DEL	182	37	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	4.05
chr10	10189277	8+0-	chr10	10202566	0+8-	DEL	13258	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.02
chr10	10220062	13+0-	chr10	10220524	0+13-	DEL	422	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	0.24
chr10	10284384	14+0-	chr10	10292025	0+14-	DEL	7629	99	14	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|14	NA
chr10	10313482	24+1-	chr10	10313837	1+25-	DEL	345	99	24	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|24	0.08
chr10	10353763	7+0-	chr10	10353850	0+7-	DEL	92	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	1.12
chr10	10363306	13+0-	chr10	10375894	0+13-	DEL	12594	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	0.00
chr10	10418939	8+0-	chr10	10421715	0+8-	DEL	2762	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.02
chr10	10504161	4+0-	chr10	10506034	0+4-	DEL	1821	80	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	NA
chr10	10533312	3+0-	chr10	10533737	0+3-	DEL	337	83	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.03
chr10	10572991	4+0-	chr10	10573070	0+4-	DEL	91	65	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.80
chr10	10631052	12+0-	chr10	10634276	0+11-	DEL	3210	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	0.01
chr10	10656503	4+0-	chr10	10657944	0+5-	DEL	1350	82	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	2.10
chr10	10660526	2+4-	chr10	10660615	2+4-	INV	-59	67	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr10	10668157	15+0-	chr10	10674626	1+15-	DEL	6444	99	14	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|14	0.01
chr10	10711025	4+11-	chr10	10711254	4+11-	INV	57	57	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr10	10711289	4+11-	chr10	10711514	0+11-	INV	94	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	0.64
chr10	10712881	22+0-	chr10	10713100	0+22-	DEL	235	99	22	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|22	NA
chr10	10715699	7+1-	chr10	10723034	0+7-	DEL	7325	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	0.00
chr10	10723737	7+0-	chr10	10724033	1+8-	DEL	282	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	0.05
chr10	10737077	5+0-	chr10	10737851	0+5-	DEL	768	84	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.04
chr10	10749863	4+0-	chr10	10750150	0+3-	DEL	239	64	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.14
chr10	10752379	17+0-	chr10	10754096	1+17-	DEL	1705	99	16	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|16	0.04
chr10	10971783	5+0-	chr10	10975347	0+5-	DEL	3480	99	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.00
chr10	10980210	6+0-	chr10	10982600	0+6-	DEL	2329	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.03
chr10	10983123	2+0-	chr10	10985839	0+2-	DEL	2627	57	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.01
chr10	11022866	2+0-	chr10	11026234	0+4-	DEL	3271	49	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.02
chr10	11026113	2+0-	chr10	11026234	0+4-	DEL	86	48	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.19
chr10	11043732	15+0-	chr10	11045047	0+15-	DEL	1299	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	0.02
chr10	11122865	18+0-	chr10	11123140	0+19-	DEL	271	99	18	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|18	0.25
chr10	11208867	9+0-	chr10	11209027	0+8-	DEL	100	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.16
chr10	11227680	11+0-	chr10	11227937	0+11-	DEL	241	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	NA
chr10	11228443	15+1-	chr10	11233851	4+18-	DEL	5407	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	0.01
chr10	11241896	17+0-	chr10	11242395	0+17-	DEL	515	99	17	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|17	NA
chr10	11266838	14+1-	chr10	11266908	0+13-	DEL	93	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	0.43
chr10	11326727	6+0-	chr10	11327014	0+6-	DEL	249	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	NA
chr10	11328981	5+0-	chr10	11335414	0+6-	DEL	6429	83	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.01
chr10	11374181	3+1-	chr10	11380982	0+5-	DEL	6775	55	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	NA
chr10	11374780	2+0-	chr10	11380982	0+5-	DEL	6168	45	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr10	11383847	10+0-	chr10	11384426	1+10-	DEL	532	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	0.02
chr10	11391837	2+0-	chr10	11392044	0+2-	DEL	111	64	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.69
chr10	11545366	7+1-	chr10	11545457	0+7-	DEL	118	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	0.36
chr10	11551440	2+0-	chr10	11551570	0+2-	DEL	84	43	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.09
chr10	11643310	19+0-	chr10	11643543	2+20-	DEL	253	99	19	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|19	NA
chr10	11676793	18+0-	chr10	11689477	0+18-	DEL	12669	99	18	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|18	0.00
chr10	11691011	3+0-	chr10	11691175	0+3-	DEL	92	69	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	2.52
chr10	11704131	4+0-	chr10	11712637	0+4-	DEL	8421	99	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.02
chr10	11763805	10+0-	chr10	11776706	0+10-	DEL	12867	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	NA
chr10	11789404	9+0-	chr10	11789654	0+9-	DEL	177	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	NA
chr10	11799541	3+0-	chr10	11799850	0+3-	DEL	251	66	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.18
chr10	11909200	6+0-	chr10	11909571	0+6-	DEL	339	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	NA
chr10	11953596	8+0-	chr10	11953787	19+10-	DEL	160	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.13
chr10	11953980	19+10-	chr10	11954289	0+18-	DEL	298	99	18	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|18	0.09
chr10	11958144	6+2-	chr10	11958272	0+6-	DEL	90	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	1.49
chr10	11960519	12+0-	chr10	11960620	0+12-	DEL	110	99	12	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|12	0.45
chr10	11986199	12+1-	chr10	11987801	2+12-	DEL	1597	99	12	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|12	0.01
chr10	11995323	12+0-	chr10	11995447	0+12-	DEL	94	99	12	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|12	0.57
chr10	11999277	8+0-	chr10	12000293	0+8-	DEL	940	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.20
chr10	12004203	15+0-	chr10	12004393	0+16-	DEL	276	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	0.07
chr10	12014977	16+0-	chr10	12015095	0+16-	DEL	112	99	16	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|16	0.50
chr10	12110226	14+1-	chr10	12111609	0+13-	DEL	1386	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	0.01
chr10	12130938	13+0-	chr10	12133889	0+14-	DEL	2920	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	0.04
chr10	12154009	9+0-	chr10	12165138	0+9-	DEL	11089	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	0.00
chr10	12177921	12+0-	chr10	12179392	0+12-	DEL	1473	99	12	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|12	NA
chr10	12187531	8+0-	chr10	12187878	0+8-	DEL	334	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.08
chr10	12190031	18+0-	chr10	12190666	0+18-	DEL	630	99	18	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|18	0.11
chr10	12192086	3+0-	chr10	12192307	0+4-	DEL	149	61	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.06
chr10	12208213	6+0-	chr10	12209365	1+7-	DEL	1172	95	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	1.00
chr10	12223591	4+0-	chr10	12250376	0+4-	DEL	26698	99	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.01
chr10	12310336	7+0-	chr10	12310532	0+7-	DEL	129	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	0.26
chr10	12314113	2+0-	chr10	12314797	0+2-	DEL	586	65	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.02
chr10	12339863	9+0-	chr10	12351180	0+9-	DEL	11279	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	1.54
chr10	12346046	8+0-	chr10	12346253	0+8-	DEL	118	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.63
chr10	12454972	4+0-	chr10	12458199	0+4-	DEL	3154	89	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.00
chr10	12599806	0+17-	chr10	12649058	0+17-	INV	49070	99	17	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|17	0.05
chr10	12671680	2+0-	chr10	12671822	2+0-	INV	-32	77	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.69
chr10	12673269	19+0-	chr10	12676423	0+18-	DEL	3161	99	18	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|18	0.02
chr10	12679623	8+0-	chr10	12683897	0+8-	DEL	4277	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	NA
chr10	12745021	14+0-	chr10	12753020	0+14-	DEL	7994	99	14	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|14	NA
chr10	12779340	2+0-	chr10	12797272	0+2-	DEL	17839	61	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	2.97
chr10	12864908	5+0-	chr10	12865153	0+5-	DEL	260	81	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.05
chr10	13034929	3+12-	chr10	13035055	0+3-	DEL	93	50	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	1.32
chr10	12867343	5+0-	chr10	12867462	0+5-	DEL	83	95	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	1.38
chr10	12949644	5+0-	chr10	12950341	0+5-	DEL	674	87	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.02
chr10	13051405	6+0-	chr10	13051672	0+6-	DEL	233	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.05
chr10	13057976	9+0-	chr10	13058133	0+9-	DEL	98	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	0.79
chr10	13065335	3+0-	chr10	13066011	0+2-	DEL	576	48	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.06
chr10	13108672	9+0-	chr10	13108926	6+6-	DEL	230	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.11
chr10	13108672	9+0-	chr10	13109195	0+9-	DEL	440	54	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.08
chr10	13109034	6+6-	chr10	13109195	0+9-	DEL	202	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.08
chr10	13127573	4+0-	chr10	13127819	0+4-	DEL	216	75	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.22
chr10	13138223	3+0-	chr10	13138512	0+3-	DEL	211	68	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.70
chr10	13282982	5+0-	chr10	13283120	0+4-	DEL	121	70	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.35
chr10	13372352	8+0-	chr10	13373535	0+8-	DEL	1166	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	NA
chr10	13403528	3+0-	chr10	13404031	0+3-	DEL	411	84	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.17
chr10	13404651	3+0-	chr10	13404839	0+3-	DEL	99	76	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.34
chr10	13451727	3+0-	chr10	13461445	0+3-	DEL	9648	69	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	NA
chr10	13535531	4+0-	chr10	13535585	4+0-	INV	-93	71	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr10	13555729	10+0-	chr10	13556436	0+10-	DEL	688	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	0.02
chr10	13665520	12+0-	chr10	13673460	0+12-	DEL	7929	99	12	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|12	0.01
chr10	13696795	23+0-	chr10	13696976	0+23-	DEL	193	99	23	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|23	NA
chr10	13699889	11+0-	chr10	13700179	0+11-	DEL	263	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	0.14
chr10	14039614	5+3-	chr10	14042790	0+4-	DEL	3120	80	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	1.76
chr10	13951194	2+0-	chr10	13951398	0+4-	DEL	143	50	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.06
chr10	13958417	16+0-	chr10	13958549	1+16-	DEL	136	99	16	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|16	0.18
chr10	14010335	3+0-	chr10	14010519	0+3-	DEL	104	75	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	1.18
chr10	14019982	7+0-	chr10	14020193	0+7-	DEL	222	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	0.31
chr10	14021237	7+0-	chr10	14023698	3+7-	DEL	2435	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	NA
chr10	14023821	3+7-	chr10	14024113	0+3-	DEL	259	64	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.05
chr10	14037563	5+0-	chr10	14038241	0+5-	DEL	594	99	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.11
chr10	14040061	6+3-	chr10	14040184	0+6-	DEL	123	91	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.19
chr10	14041101	7+0-	chr10	14041314	0+7-	DEL	154	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	0.37
chr10	14042302	24+3-	chr10	14042545	0+22-	DEL	248	99	22	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|22	0.05
chr10	14046528	4+0-	chr10	14054514	1+4-	DEL	7915	95	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.02
chr10	14065394	6+1-	chr10	14065648	27+7-	DEL	246	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	NA
chr10	14065840	27+7-	chr10	14066122	2+27-	DEL	290	99	27	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|27	0.10
chr10	14071646	15+0-	chr10	14071992	0+15-	DEL	335	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	0.08
chr10	14073268	3+0-	chr10	14073681	0+3-	DEL	379	57	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.03
chr10	14076552	15+0-	chr10	14085825	0+15-	DEL	9282	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	0.00
chr10	14111731	11+0-	chr10	14115774	0+11-	DEL	4009	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	0.01
chr10	14173173	14+0-	chr10	14173987	0+14-	DEL	824	99	14	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|14	NA
chr10	14184965	8+0-	chr10	14191478	0+7-	DEL	6455	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	0.01
chr10	14195658	24+1-	chr10	14202002	0+23-	DEL	6350	99	23	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|23	0.00
chr10	14208177	4+0-	chr10	14208284	0+4-	DEL	95	68	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.11
chr10	14210375	22+0-	chr10	14213927	0+22-	DEL	3565	99	22	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|22	NA
chr10	14215450	17+0-	chr10	14215698	0+17-	DEL	267	99	17	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|17	NA
chr10	14223193	4+0-	chr10	14224001	0+4-	DEL	710	99	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	NA
chr10	14237269	12+0-	chr10	14253724	0+12-	DEL	16461	99	12	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|12	NA
chr10	14278505	4+0-	chr10	14281869	0+4-	DEL	3288	89	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	NA
chr10	14349119	7+1-	chr10	14349219	7+1-	INV	-104	91	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	NA
chr10	14365295	25+0-	chr10	14370080	0+25-	DEL	4789	99	25	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|25	0.00
chr10	14415392	4+0-	chr10	14415490	0+4-	DEL	81	71	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	1.26
chr10	14457351	5+0-	chr10	14457465	0+5-	DEL	108	83	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	1.22
chr10	14562286	18+0-	chr10	14562537	0+18-	DEL	226	99	18	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|18	0.42
chr10	14578029	23+0-	chr10	14578343	1+24-	DEL	315	99	23	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|23	0.13
chr10	14583870	10+1-	chr10	14584184	1+10-	DEL	337	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	NA
chr10	14585402	4+0-	chr10	14585548	0+4-	DEL	90	82	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	1.01
chr10	14676997	17+0-	chr10	14677465	0+18-	DEL	456	99	17	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|17	NA
chr10	14708464	3+0-	chr10	14708789	0+3-	DEL	245	74	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.13
chr10	14716630	3+3-	chr10	14716964	3+3-	DEL	81	42	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	NA
chr10	14724146	3+0-	chr10	14724311	0+3-	DEL	98	66	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	1.90
chr10	14725116	15+0-	chr10	14731187	0+15-	DEL	6047	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	3.44
chr10	14748774	21+2-	chr10	14748981	0+21-	DEL	268	99	21	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|21	0.06
chr10	14797103	22+0-	chr10	14797621	0+22-	DEL	526	99	22	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|22	0.03
chr10	14930364	23+6-	chr10	14938155	0+22-	DEL	7912	99	21	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|21	NA
chr10	14820359	5+1-	chr10	14820551	0+4-	DEL	121	79	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.13
chr10	14872237	3+0-	chr10	14874075	0+3-	DEL	1765	65	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.02
chr10	14882311	10+0-	chr10	14882502	0+8-	DEL	134	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	0.27
chr10	14882311	10+0-	chr10	14894547	1+3-	DEL	12244	62	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.08
chr10	14915962	9+0-	chr10	14916182	0+9-	DEL	156	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	0.06
chr10	14950267	7+0-	chr10	14950408	1+8-	DEL	86	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	1.04
chr10	14989570	11+0-	chr10	15002965	0+12-	DEL	13353	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	0.00
chr10	15050412	12+0-	chr10	15051031	0+12-	DEL	623	99	12	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|12	0.07
chr10	15111593	4+0-	chr10	15111937	0+4-	DEL	246	99	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.12
chr10	15123269	7+0-	chr10	15123924	0+7-	DEL	610	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	0.09
chr10	15126010	16+0-	chr10	15126334	0+16-	DEL	332	99	16	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|16	0.04
chr10	15128869	15+0-	chr10	15137127	0+16-	DEL	8263	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	NA
chr10	15168228	19+1-	chr10	15168568	0+18-	DEL	343	99	18	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|18	0.20
chr10	15169268	19+0-	chr10	15169606	0+19-	DEL	347	99	19	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|19	0.04
chr10	15170961	5+0-	chr10	15171485	0+5-	DEL	471	98	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.03
chr10	15171865	12+0-	chr10	15172293	0+13-	DEL	401	99	12	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|12	0.03
chr10	15188667	18+1-	chr10	15188921	0+13-	DEL	250	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	0.11
chr10	15189779	6+0-	chr10	15189978	0+6-	DEL	172	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.26
chr10	15195359	7+0-	chr10	15198951	1+7-	DEL	3550	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	0.00
chr10	15201464	4+0-	chr10	15204943	0+4-	DEL	3414	80	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.00
chr10	15217867	4+0-	chr10	15218107	0+4-	DEL	247	67	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.06
chr10	15308352	6+0-	chr10	15308535	0+6-	DEL	108	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.56
chr10	15310050	14+0-	chr10	15323230	1+13-	DEL	13211	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	NA
chr10	15347245	5+0-	chr10	15347334	0+5-	DEL	93	82	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.61
chr10	15385635	4+0-	chr10	15391238	0+3-	DEL	5508	68	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.02
chr10	15403687	13+1-	chr10	15403799	0+13-	DEL	101	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	0.52
chr10	15415037	22+4-	chr10	15415336	22+4-	INV	-30	54	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr10	15415371	22+4-	chr10	15419540	1+22-	DEL	4215	99	22	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|22	0.01
chr10	15440802	2+0-	chr10	15441940	0+3-	DEL	1067	49	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.04
chr10	15453755	6+1-	chr10	15522683	0+6-	DEL	68838	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	1.10
chr10	15461506	5+1-	chr10	15461580	0+5-	DEL	90	81	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.84
chr10	15504899	2+0-	chr10	15505071	2+0-	INV	-2	71	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	1.54
chr10	15549298	4+0-	chr10	15549506	0+4-	DEL	170	77	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	NA
chr10	15550979	2+0-	chr10	15557485	0+2-	DEL	6436	49	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.01
chr10	15572595	2+0-	chr10	15572769	2+0-	INV	-17	73	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	1.82
chr10	15687293	8+2-	chr10	15687426	8+2-	INV	-41	87	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	NA
chr10	15702533	9+0-	chr10	15707648	0+3-	DEL	5042	64	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	NA
chr10	15743819	3+0-	chr10	15743911	0+3-	DEL	84	52	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	1.79
chr10	15767796	5+0-	chr10	15772548	0+11-	DEL	4679	65	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.01
chr10	15769543	7+2-	chr10	15772548	0+11-	DEL	2993	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	NA
chr10	15802667	3+5-	chr10	15802995	3+5-	DEL	87	42	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	NA
chr10	15848519	2+0-	chr10	15848956	0+2-	DEL	369	48	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr10	15854317	12+1-	chr10	15854578	5+11-	DEL	261	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	0.31
chr10	15854742	5+11-	chr10	15855372	0+5-	DEL	610	90	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.07
chr10	15877301	19+0-	chr10	15877567	0+19-	DEL	247	99	19	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|19	0.15
chr10	15882157	10+0-	chr10	15884987	1+11-	DEL	2798	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	0.06
chr10	15890783	2+2-	chr10	15890928	2+2-	INV	-81	62	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr10	15917788	6+0-	chr10	15918155	0+6-	DEL	317	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	NA
chr10	15939853	7+0-	chr10	15940072	0+7-	DEL	128	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	0.06
chr10	15941135	5+0-	chr10	15941567	0+5-	DEL	344	99	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.10
chr10	15951166	8+2-	chr10	15951429	9+8-	DEL	224	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	NA
chr10	15951552	9+8-	chr10	15952528	0+8-	DEL	962	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	NA
chr10	15968838	2+0-	chr10	15971092	8+2-	DEL	2167	51	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr10	15976462	7+0-	chr10	15983440	22+8-	DEL	7130	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	NA
chr10	16261260	5+0-	chr10	16262574	1+7-	DEL	1297	74	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	NA
chr10	14647441	2+0-	chr10	16085305	6+3-	INV	1437603	60	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	1.61
chr10	15971184	8+2-	chr10	15971488	1+8-	DEL	259	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.04
chr10	15975206	10+0-	chr10	15975662	0+10-	DEL	457	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	0.12
chr10	15984994	5+0-	chr10	15985630	0+5-	DEL	613	90	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	NA
chr10	15992012	11+0-	chr10	15992196	4+7-	DEL	165	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	0.14
chr10	15992012	11+0-	chr10	15992513	0+8-	DEL	425	67	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.09
chr10	15992258	4+7-	chr10	15992513	0+8-	DEL	233	76	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	NA
chr10	15999008	2+0-	chr10	15999133	0+2-	DEL	84	42	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	1.52
chr10	16003379	6+0-	chr10	16003629	0+6-	DEL	155	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.16
chr10	16148582	2+0-	chr10	16148790	0+3-	DEL	160	43	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	5.75
chr10	16214048	23+0-	chr10	16217994	2+23-	DEL	3911	99	23	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|23	NA
chr10	16274764	13+2-	chr10	16275043	14+12-	DEL	257	99	12	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|12	0.05
chr10	16275167	14+12-	chr10	16275426	0+14-	DEL	245	99	14	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|14	0.16
chr10	16276577	14+0-	chr10	16276748	0+14-	DEL	156	99	14	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|14	0.15
chr10	16282628	4+0-	chr10	16282950	0+4-	DEL	227	99	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.09
chr10	16293410	16+1-	chr10	16293614	0+16-	DEL	207	99	16	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|16	0.06
chr10	16312533	16+0-	chr10	16313740	0+16-	DEL	1220	99	16	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|16	0.01
chr10	16328472	2+0-	chr10	16328574	1+2-	DEL	80	42	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	1.11
chr10	16460895	21+0-	chr10	16473886	0+21-	DEL	12987	99	21	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|21	0.00
chr10	16484126	5+0-	chr10	16485239	0+5-	DEL	1113	86	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.01
chr10	16489200	4+0-	chr10	16489443	0+7-	DEL	245	79	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	NA
chr10	16492574	20+0-	chr10	16492717	0+20-	DEL	139	99	20	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|20	0.17
chr10	16499179	3+1-	chr10	16499731	0+3-	DEL	504	52	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	NA
chr10	16535090	1+5-	chr10	16535236	1+5-	INV	-1	62	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr10	16606618	3+0-	chr10	16606957	0+3-	DEL	249	79	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.04
chr10	16610176	15+0-	chr10	16610322	1+15-	DEL	132	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	NA
chr10	16620436	15+0-	chr10	16620712	0+16-	DEL	254	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	0.15
chr10	16637971	6+0-	chr10	16638199	0+6-	DEL	147	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.06
chr10	16644385	9+0-	chr10	16644708	0+9-	DEL	275	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	0.21
chr10	16674246	0+2-	chr10	16675371	0+2-	INV	934	81	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	1.51
chr10	16710650	4+0-	chr10	16710682	4+0-	INV	-115	75	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr10	16744127	24+0-	chr10	16749886	0+23-	DEL	5756	99	23	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|23	0.01
chr10	16824915	17+0-	chr10	16825084	0+17-	DEL	168	99	17	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|17	0.45
chr10	16855815	15+0-	chr10	16860911	0+15-	DEL	5074	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	0.01
chr10	16866755	13+1-	chr10	16866873	13+1-	INV	-29	64	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr10	16866908	13+1-	chr10	16867042	0+10-	DEL	126	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	0.09
chr10	16872131	14+0-	chr10	16884053	0+14-	DEL	11933	99	14	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|14	NA
chr10	16887032	4+0-	chr10	16890678	0+4-	DEL	3623	74	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.00
chr10	17055231	3+0-	chr10	17063040	0+3-	DEL	7735	68	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.01
chr10	17146045	4+0-	chr10	17146601	0+4-	DEL	505	78	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.13
chr10	17275150	4+0-	chr10	17275463	0+4-	DEL	223	99	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.61
chr10	17311345	4+1-	chr10	17311537	0+4-	DEL	131	77	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.13
chr10	17322596	15+0-	chr10	17323398	0+15-	DEL	778	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	0.05
chr10	17373075	15+1-	chr10	17373332	0+9-	DEL	252	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	0.05
chr10	17376640	15+0-	chr10	17376996	0+15-	DEL	353	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	0.16
chr10	17381331	5+0-	chr10	17381499	0+5-	DEL	87	99	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.60
chr10	17383498	11+0-	chr10	17385028	0+12-	DEL	1522	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	0.05
chr10	17422044	10+0-	chr10	17431095	0+10-	DEL	9053	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	0.00
chr10	17491315	10+0-	chr10	17492592	0+10-	DEL	1241	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	0.02
chr10	14066472	2+2-	chr10	17496703	0+2-	INV	3430044	79	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	1.76
chr10	17498971	12+1-	chr10	17499047	0+10-	DEL	136	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	0.14
chr10	17624152	2+0-	chr10	17636872	1+3-	DEL	12670	51	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.00
chr10	17639225	8+1-	chr10	17642452	0+9-	DEL	3179	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.01
chr10	17719161	7+3-	chr10	17719323	0+3-	DEL	96	44	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.93
chr10	17816532	6+0-	chr10	17816762	0+6-	DEL	217	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.06
chr10	17819484	10+0-	chr10	17830830	0+10-	DEL	11308	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	0.01
chr10	18176894	1+7-	chr10	18178640	1+3-	INV	1564	89	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.34
chr10	17854924	3+0-	chr10	17855154	0+3-	DEL	140	83	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.52
chr10	17898268	16+0-	chr10	17898631	13+11-	DEL	367	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	0.04
chr10	17898268	16+0-	chr10	17899053	0+18-	DEL	703	79	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.02
chr10	17898714	13+11-	chr10	17899053	0+18-	DEL	350	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	NA
chr10	17902775	11+0-	chr10	17902907	0+12-	DEL	107	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	0.36
chr10	17930927	5+0-	chr10	17930992	5+0-	INV	-82	70	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr10	18031592	14+0-	chr10	18031934	0+14-	DEL	349	99	14	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|14	NA
chr10	18038164	8+0-	chr10	18038294	8+0-	INV	-75	99	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	NA
chr10	18124525	10+0-	chr10	18125247	0+10-	DEL	697	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	0.08
chr10	18149916	19+0-	chr10	18150159	0+19-	DEL	250	99	19	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|19	0.05
chr10	18220660	10+0-	chr10	18220800	1+11-	DEL	118	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	0.17
chr10	18231226	32+0-	chr10	18231325	0+32-	DEL	106	99	32	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|32	0.68
chr10	18289864	21+0-	chr10	18294317	0+21-	DEL	4436	99	21	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|21	0.01
chr10	18297410	14+2-	chr10	18297709	0+11-	DEL	280	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	0.18
chr10	18340405	0+4-	chr10	18340428	0+4-	INV	-125	77	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr10	18388277	2+2-	chr10	18388467	2+2-	INV	-119	59	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr10	18529750	5+1-	chr10	18530035	5+1-	INV	-48	55	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr10	18571165	8+0-	chr10	18571559	0+8-	DEL	392	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	NA
chr10	18606211	6+13-	chr10	18620599	8+14-	DEL	14766	49	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	3.84
chr10	18600705	9+0-	chr10	18620599	8+14-	DEL	20077	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	2.80
chr10	18572342	12+0-	chr10	18572447	0+11-	DEL	89	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	1.19
chr10	18619297	12+0-	chr10	18619372	0+12-	DEL	97	99	12	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|12	0.28
chr10	18621474	2+0-	chr10	18627977	1+2-	DEL	6403	55	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.01
chr10	18655621	4+0-	chr10	18655842	0+4-	DEL	146	95	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.24
chr10	18690005	4+1-	chr10	18690060	4+1-	INV	-92	71	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr10	18711398	4+0-	chr10	18712396	1+4-	DEL	919	81	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.01
chr10	18713066	3+0-	chr10	18714223	0+3-	DEL	1087	71	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.14
chr10	18724172	8+0-	chr10	18724362	0+8-	DEL	184	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.07
chr10	18765785	17+0-	chr10	18765895	0+15-	DEL	112	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	0.10
chr10	18775724	2+3-	chr10	18775961	2+3-	INV	-28	57	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr10	18779451	22+1-	chr10	18779758	1+23-	DEL	341	99	22	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|22	NA
chr10	18780200	2+5-	chr10	18780342	2+5-	INV	-137	62	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr10	18720125	3+0-	chr10	18953889	1+6-	DEL	233759	60	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	2.58
chr10	18938492	3+5-	chr10	18953889	1+6-	DEL	15308	62	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	1.10
chr10	18921517	4+0-	chr10	18934166	0+3-	DEL	12658	57	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.08
chr10	18991563	12+0-	chr10	18992189	1+12-	DEL	619	99	12	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|12	0.09
chr10	18993149	21+0-	chr10	18993501	0+24-	DEL	345	99	20	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|20	0.12
chr10	18997387	13+0-	chr10	18998395	2+13-	DEL	1019	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	NA
chr10	19008262	19+0-	chr10	19008761	0+19-	DEL	506	99	19	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|19	0.03
chr10	19027956	2+0-	chr10	19028120	0+2-	DEL	98	47	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.84
chr10	19034601	6+0-	chr10	19034676	0+6-	DEL	87	98	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	1.52
chr10	19042153	9+1-	chr10	19042628	0+9-	DEL	457	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	0.27
chr10	19049777	4+0-	chr10	19050172	1+4-	DEL	319	90	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.21
chr10	19086824	3+0-	chr10	19086992	0+3-	DEL	86	75	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	2.24
chr10	19104456	7+0-	chr10	19104633	0+7-	DEL	141	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	0.07
chr10	19122188	8+0-	chr10	19122396	1+8-	DEL	248	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	NA
chr10	19123568	2+0-	chr10	19123723	1+3-	DEL	90	47	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	1.52
chr10	19144457	7+1-	chr10	19144605	0+7-	DEL	101	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	0.42
chr10	19174902	9+2-	chr10	19176407	0+9-	DEL	1452	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	0.18
chr10	19176909	15+0-	chr10	19189946	0+15-	DEL	13045	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	0.00
chr10	19223959	6+0-	chr10	19224053	0+6-	DEL	94	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	1.41
chr10	19234887	15+0-	chr10	19235038	0+15-	DEL	116	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	0.25
chr10	19242075	5+0-	chr10	19243953	0+5-	DEL	1860	90	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.02
chr10	19340156	9+0-	chr10	19340802	0+9-	DEL	578	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	0.02
chr10	19376421	10+0-	chr10	19376786	0+10-	DEL	337	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	0.08
chr10	19377725	3+0-	chr10	19377837	0+3-	DEL	81	57	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	1.65
chr10	19381765	15+0-	chr10	19382486	0+15-	DEL	701	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	0.02
chr10	19386573	9+0-	chr10	19387809	0+9-	DEL	1182	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	0.04
chr10	19398565	15+0-	chr10	19398859	0+15-	DEL	296	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	NA
chr10	19416191	5+0-	chr10	19416397	0+5-	DEL	133	99	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.19
chr10	19432326	19+0-	chr10	19432779	0+19-	DEL	450	99	19	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|19	0.06
chr10	19440720	7+1-	chr10	19448572	1+7-	DEL	7877	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	0.01
chr10	19472112	13+0-	chr10	19472453	0+13-	DEL	338	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	0.04
chr10	19486297	15+0-	chr10	19501759	0+15-	DEL	15462	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	0.00
chr10	19504480	6+0-	chr10	19510964	0+6-	DEL	6412	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.01
chr10	19519191	3+0-	chr10	19519379	1+2-	DEL	92	46	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	3.41
chr10	19553166	15+0-	chr10	19553419	0+15-	DEL	252	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	0.05
chr10	19605518	8+0-	chr10	19605879	0+8-	DEL	334	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.15
chr10	19654807	4+0-	chr10	19654952	2+2-	DEL	108	48	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.17
chr10	19654807	4+0-	chr10	19661448	0+4-	DEL	6548	39	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.01
chr10	19655029	2+2-	chr10	19661448	0+4-	DEL	6435	39	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr10	19699671	5+0-	chr10	19703340	0+5-	DEL	3583	99	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.01
chr10	19720635	20+0-	chr10	19720959	0+20-	DEL	327	99	20	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|20	NA
chr10	19731267	17+0-	chr10	19731809	1+18-	DEL	523	99	17	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|17	0.11
chr10	19824040	8+0-	chr10	19824297	0+8-	DEL	196	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	NA
chr10	19829976	3+0-	chr10	19831658	0+3-	DEL	1660	54	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	NA
chr10	19844445	3+0-	chr10	19847022	0+3-	DEL	2499	71	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.01
chr10	19848711	8+0-	chr10	19849015	0+8-	DEL	236	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.09
chr10	19851723	22+0-	chr10	19853552	17+22-	DEL	1841	99	22	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|22	0.02
chr10	19853787	17+22-	chr10	19855994	1+17-	DEL	2206	99	17	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|17	0.02
chr10	19866415	17+0-	chr10	19867091	18+17-	DEL	695	99	17	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|17	NA
chr10	19867285	18+17-	chr10	19868821	0+19-	DEL	1551	99	18	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|18	NA
chr10	19880059	14+0-	chr10	19880309	1+14-	DEL	222	99	14	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|14	0.05
chr10	19906006	3+0-	chr10	19906136	0+3-	DEL	85	61	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	3.04
chr10	19926568	15+0-	chr10	19926680	0+15-	DEL	102	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	1.14
chr10	19927696	11+1-	chr10	19927828	0+11-	DEL	127	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	0.09
chr10	19944538	9+0-	chr10	19944984	0+9-	DEL	423	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	0.06
chr10	19959960	6+0-	chr10	19960058	0+6-	DEL	103	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.23
chr10	20009038	20+0-	chr10	20010044	0+20-	DEL	1009	99	20	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|20	0.04
chr10	20014236	18+1-	chr10	20016647	1+18-	DEL	2432	99	17	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|17	0.01
chr10	20044409	0+4-	chr10	20044467	0+4-	INV	-89	71	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr10	20049558	9+0-	chr10	20056025	1+10-	DEL	6422	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	0.02
chr10	20103906	4+0-	chr10	20107979	0+4-	DEL	3983	97	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.06
chr10	20122369	17+0-	chr10	20122658	0+17-	DEL	268	99	17	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|17	0.19
chr10	20162741	3+0-	chr10	20163143	0+3-	DEL	362	60	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	NA
chr10	20205662	8+0-	chr10	20206028	0+8-	DEL	352	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.11
chr10	20212944	5+1-	chr10	20213129	0+4-	DEL	128	71	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.21
chr10	20215140	11+0-	chr10	20216235	0+11-	DEL	1087	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	0.03
chr10	20248956	21+0-	chr10	20249193	0+21-	DEL	231	99	21	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|21	0.22
chr10	20286609	7+0-	chr10	20286892	0+7-	DEL	192	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	0.05
chr10	20294908	7+0-	chr10	20295137	0+7-	DEL	165	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	NA
chr10	20296878	3+0-	chr10	20297147	0+3-	DEL	173	80	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	2.95
chr10	20300261	7+0-	chr10	20300559	0+7-	DEL	248	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	NA
chr10	20308998	6+0-	chr10	20309213	0+6-	DEL	132	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.06
chr10	18919858	6+6-	chr10	20396696	0+3-	DEL	1476873	49	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	2.33
chr10	20313480	7+0-	chr10	20314634	0+7-	DEL	1161	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	NA
chr10	20319953	3+0-	chr10	20326365	0+3-	DEL	6324	77	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.74
chr10	20327190	10+0-	chr10	20327496	0+10-	DEL	248	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	0.18
chr10	20352569	5+0-	chr10	20352749	2+5-	DEL	133	94	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.71
chr10	20384317	2+6-	chr10	20384390	2+6-	INV	-99	69	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr10	20492821	5+3-	chr10	20493254	0+5-	DEL	404	95	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.13
chr10	20495410	8+0-	chr10	20495841	0+8-	DEL	347	99	8	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|8	0.03
chr10	20541763	12+4-	chr10	20541983	12+4-	INV	-81	58	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr10	20542018	12+4-	chr10	20550159	0+12-	DEL	8117	99	12	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|12	0.01
chr10	20577421	23+0-	chr10	20589044	1+23-	DEL	11632	99	23	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|23	0.00
chr10	20630082	24+0-	chr10	20630389	0+24-	DEL	312	99	24	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|24	0.22
chr10	20709705	5+0-	chr10	20709865	0+5-	DEL	92	99	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	2.18
chr10	20836851	24+29-	chr10	20861824	25+28-	INV	24250	99	52	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|52	3.17
chr10	20878822	6+0-	chr10	20878952	1+6-	DEL	115	95	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.18
chr10	20949712	3+0-	chr10	20953711	0+4-	DEL	3906	71	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.02
chr10	20956478	5+11-	chr10	20971110	0+5-	DEL	14617	77	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	1.33
chr10	20973704	6+0-	chr10	20977791	0+6-	DEL	3994	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	0.00
chr10	20984336	7+0-	chr10	20984861	0+7-	DEL	450	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	NA
chr10	21005796	25+0-	chr10	21005942	1+26-	DEL	153	99	25	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|25	NA
chr10	21018741	3+0-	chr10	21018921	0+3-	DEL	83	87	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	2.83
chr10	21061679	16+0-	chr10	21073387	0+16-	DEL	11696	99	16	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|16	NA
chr10	21080804	21+10-	chr10	21083906	0+15-	DEL	3083	99	15	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|15	0.01
chr10	21118204	6+3-	chr10	21122903	0+6-	DEL	4745	99	6	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|6	NA
chr10	21131312	10+0-	chr10	21132300	0+10-	DEL	937	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	0.18
chr10	21205460	3+0-	chr10	21219386	0+3-	DEL	13843	69	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.04
chr10	21230086	4+0-	chr10	21230127	4+0-	INV	-106	73	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr10	21265297	13+0-	chr10	21265420	0+13-	DEL	106	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	0.48
chr10	21267326	5+0-	chr10	21267513	0+5-	DEL	99	99	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.89
chr10	21368077	5+0-	chr10	21368155	0+5-	DEL	89	82	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.27
chr10	21394405	4+0-	chr10	21394603	0+4-	DEL	103	99	4	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|4	0.20
chr10	21459222	2+1-	chr10	21459364	1+2-	DEL	97	47	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	4.72
chr10	21493387	15+1-	chr10	21504692	0+14-	DEL	11325	99	14	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|14	0.00
chr10	21527204	20+0-	chr10	21531190	0+20-	DEL	3994	99	20	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|20	NA
chr10	21554070	16+0-	chr10	21557857	0+16-	DEL	3813	99	16	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|16	0.01
chr10	21595440	4+1-	chr10	21595748	1+4-	DEL	308	37	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	5.31
chr10	21597901	19+0-	chr10	21598065	0+19-	DEL	140	99	19	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|19	0.15
chr10	21672548	11+0-	chr10	21673136	13+11-	DEL	592	99	11	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|11	0.05
chr10	21673349	13+11-	chr10	21673658	0+13-	DEL	309	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	NA
chr10	21684982	5+0-	chr10	21689548	0+5-	DEL	4500	99	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.02
chr10	21716384	18+0-	chr10	21716837	0+18-	DEL	440	99	18	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|18	0.12
chr10	21746240	16+0-	chr10	21746491	0+16-	DEL	246	99	16	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|16	0.21
chr10	21767847	19+0-	chr10	21767949	2+19-	DEL	95	99	18	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|18	0.67
chr10	21792882	14+0-	chr10	21793770	0+14-	DEL	887	99	14	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|14	0.02
chr10	21821158	3+0-	chr10	21822225	0+3-	DEL	993	66	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	0.04
chr10	21842004	16+0-	chr10	21842790	0+16-	DEL	788	99	16	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|16	0.02
chr10	21917163	9+0-	chr10	21921896	0+9-	DEL	4734	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	0.01
chr10	22183626	13+5-	chr10	22184632	0+13-	DEL	1097	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	0.03
chr10	22025792	8+1-	chr10	22025912	0+7-	DEL	92	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	1.37
chr10	22038876	2+0-	chr10	22039048	0+2-	DEL	95	51	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	1.98
chr10	22068614	19+0-	chr10	22069732	3+22-	DEL	1114	99	19	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|19	0.04
chr10	22143427	8+3-	chr10	22143702	0+5-	DEL	261	87	5	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|5	0.05
chr10	22178030	13+0-	chr10	22178278	0+13-	DEL	243	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	0.05
chr10	22300477	21+1-	chr10	22306183	0+21-	DEL	5714	99	21	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|21	NA
chr10	22330002	13+0-	chr10	22330290	0+13-	DEL	269	99	13	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|13	NA
chr10	22588217	16+11-	chr10	22591334	15+16-	DEL	3437	99	16	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|16	1.16
chr10	15253742	20+0-	chr10	22517096	0+3-	DEL	7263284	64	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	2.30
chr10	19419238	0+3-	chr10	22600434	0+5-	INV	3181001	91	3	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|3	2.53
chr10	22369095	10+0-	chr10	22369462	0+10-	DEL	347	99	10	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|10	0.08
chr10	22372359	7+0-	chr10	22372814	0+7-	DEL	434	99	7	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|7	NA
chr10	22402722	12+0-	chr10	22408475	0+12-	DEL	5750	99	12	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|12	NA
chr10	22439411	16+0-	chr10	22440822	0+16-	DEL	1396	99	16	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|16	0.04
chr10	22444822	2+0-	chr10	22449343	0+2-	DEL	4437	55	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	0.03
chr10	22505649	0+4-	chr10	22505654	0+4-	INV	-143	81	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	NA
chr10	22522763	9+0-	chr10	22522874	0+9-	DEL	96	99	9	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|9	0.52
chr10	22678621	34+0-	chr10	22679240	0+32-	DEL	629	99	32	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|32	0.46
chr10	22777683	2+0-	chr10	22777832	0+2-	DEL	91	45	2	/public07/yaowen/intansv/zs97_ncgr/ZS97.bam|2	4.21
